magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l34d0 >>
<< l21d0 >>
<< l36d0 >>
<< l32d0 >>
<< labels >>
rlabel l34d10 -0.388 -0.1735 -0.388 -0.1735 0 out
rlabel l34d10 -0.516 -0.189 -0.516 -0.189 0 in1
rlabel l34d10 -0.1145 -0.1715 -0.1145 -0.1715 0 in2
rlabel l34d10 0.0155 -0.171 0.0155 -0.171 0 cntrl
rlabel l34d10 -0.3665 0.108 -0.3665 0.108 0 vdd
rlabel l34d10 -0.3575 -0.4165 -0.3575 -0.4165 0 vss
use pfetx2414 pfetx2414_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2419 nfetx2419_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_3
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_4
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_5
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_6
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2419 nfetx2419_2
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use via_devx2431 via_devx2431_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2431 via_devx2431_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use pfetx2414 pfetx2414_2
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_7
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_8
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_9
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_10
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2419 nfetx2419_3
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use via_devx2431 via_devx2431_3
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx2431 via_devx2431_4
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use pfetx2414 pfetx2414_3
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_11
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2430 via_devx2430_12
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
<< end >>
