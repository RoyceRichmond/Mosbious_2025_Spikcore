* NGSPICE file created from DFF_10_row.ext - technology: gf180mcuD

.subckt DFF_10_row_pex D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8]
+ gc[9] gc[10] PHI_1 PHI_2 EN VDD VSS
X0 a_20582_38# a_20238_158# VSS.t62 VSS.t61 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X1 a_29738_n384# a_29270_n402# VDD.t282 VDD.t281 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 a_32570_n387# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t166 VSS.t165 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X3 VSS.t325 a_1862_38# a_1762_n387# VSS.t324 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X4 a_8102_38# a_7758_158# VSS.t176 VSS.t175 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X5 VDD.t62 a_20238_158# Q[4].t1 VDD.t61 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X6 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t0 a_27943_n425# VSS.t224 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X7 a_55214_158# a_54230_n402# a_55066_158# VDD.t203 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X8 a_5538_n387# a_4310_n402# a_5294_158# VSS.t153 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X9 VDD.t26 a_14342_38# a_14202_158# VDD.t25 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X10 VSS.t108 a_36838_38# a_36738_n387# VSS.t107 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X11 VSS.t243 PHI_1.t0 a_29270_n402# VSS.t242 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X12 a_29738_n384# a_29270_n402# VSS.t274 VSS.t273 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X13 VSS.t158 a_30254_158# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t157 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X14 VSS.t217 PHI_2.t0 a_534_n402# VSS.t216 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X15 VDD.t100 a_49318_38# a_49178_158# VDD.t99 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X16 a_11738_158# a_11018_n384# a_11534_158# VDD.t267 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X17 a_23866_158# Q[4].t2 VDD.t141 VDD.t140 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X18 VSS.t263 a_32718_158# Q[6].t0 VSS.t262 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X19 VSS.t197 a_45542_38# a_45442_n387# VSS.t196 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X20 gc[2].t1 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t106 VDD.t105 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X21 gc[2].t0 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t112 VSS.t111 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X22 a_21703_n425# Q[4].t3 VSS.t240 VSS.t239 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X23 a_38958_158# a_37974_n402# a_38810_158# VDD.t54 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X24 VSS.t219 PHI_2.t1 a_37974_n402# VSS.t218 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X25 a_38442_n384# a_37974_n402# VSS.t54 VSS.t53 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X26 VSS.t6 a_11878_38# a_11778_n387# VSS.t5 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X27 a_45198_158# a_44214_n402# a_45050_158# VDD.t24 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X28 a_42734_158# a_42218_n384# a_42586_n387# VSS.t241 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X29 a_49218_n387# a_47990_n402# a_48974_158# VSS.t9 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X30 a_55558_38# a_55214_158# VDD.t151 VDD.t150 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X31 VSS.t245 PHI_1.t1 a_41750_n402# VSS.t244 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X32 a_55558_38# a_55214_158# VSS.t147 VSS.t146 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X33 gc[8].t0 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t307 VSS.t306 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X34 VDD.t251 PHI_1.t2 a_10550_n402# VDD.t250 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X35 a_11878_38# a_11534_158# VDD.t339 VDD.t338 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X36 a_13482_n384# a_13014_n402# VDD.t57 VDD.t56 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X37 VSS.t114 a_20582_38# a_20482_n387# VSS.t113 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X38 VDD.t33 a_n946_158# DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t32 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X39 a_26822_38# a_26478_158# VSS.t139 VSS.t138 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X40 VSS.t234 a_8102_38# a_8002_n387# VSS.t233 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X41 VSS.t116 PHI_2.t2 a_13014_n402# VSS.t115 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X42 a_24258_n387# a_23030_n402# a_24014_158# VSS.t284 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X43 a_55418_158# a_54698_n384# a_55214_158# VDD.t0 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X44 a_50922_n384# a_50454_n402# VSS.t46 VSS.t45 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X45 VSS.t118 PHI_2.t3 a_50454_n402# VSS.t117 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X46 a_n1094_n387# D_in.t0 VSS.t289 VSS.t288 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X47 VDD.t180 a_7758_158# Q[2].t1 VDD.t179 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X48 a_32718_158# a_31734_n402# a_32570_158# VDD.t43 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X49 a_42586_n387# Q[7].t2 VSS.t185 VSS.t184 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X50 VDD.t116 PHI_2.t4 a_56694_n402# VDD.t115 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X51 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t1 a_21703_n425# VSS.t225 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X52 a_26822_38# a_26478_158# VDD.t137 VDD.t136 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X53 a_7758_158# a_7242_n384# a_7610_n387# VSS.t128 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X54 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t2 a_9223_n425# VSS.t226 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X55 a_26722_n387# a_25494_n402# a_26478_158# VSS.t150 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X56 VDD.t110 PHI_2.t5 a_13014_n402# VDD.t109 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X57 gc[5].t0 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t183 VSS.t182 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X58 a_57162_n384# a_56694_n402# VDD.t220 VDD.t219 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X59 VSS.t271 a_18118_38# a_18018_n387# VSS.t270 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X60 VDD.t108 a_20582_38# a_20442_158# VDD.t107 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X61 a_51290_n387# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t64 VSS.t63 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X62 a_45050_n387# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t266 VSS.t265 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X63 VDD.t236 EN.t3 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t235 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X64 VSS.t320 a_55558_38# a_55458_n387# VSS.t319 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X65 VDD.t224 a_48974_158# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t223 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X66 a_1002_n384# a_534_n402# VDD.t67 VDD.t66 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X67 a_7242_n384# a_6774_n402# VDD.t215 VDD.t214 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X68 a_5146_n387# Q[1].t2 VSS.t228 VSS.t227 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X69 VDD.t332 a_55558_38# a_55418_158# VDD.t331 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X70 a_48458_n384# a_47990_n402# VSS.t8 VSS.t7 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X71 VSS.t230 PHI_1.t3 a_47990_n402# VSS.t229 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X72 VSS.t301 a_42734_158# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t300 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X73 a_n946_158# a_n1462_n384# a_n1094_n387# VSS.t58 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X74 a_32922_158# a_32202_n384# a_32718_158# VDD.t266 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X75 a_45050_158# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t274 VDD.t273 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X76 VDD.t238 EN.t4 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t237 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X77 a_51290_158# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t64 VDD.t63 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X78 VDD.t228 PHI_1.t4 a_47990_n402# VDD.t227 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X79 a_1862_38# a_1518_158# VSS.t13 VSS.t12 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X80 gc[7].t0 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t87 VSS.t86 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X81 gc[8].t1 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t311 VDD.t310 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X82 a_24218_158# a_23498_n384# a_24014_158# VDD.t38 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X83 a_36346_158# Q[6].t2 VDD.t320 VDD.t319 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X84 a_57162_n384# a_56694_n402# VSS.t215 VSS.t214 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X85 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[1].t3 VDD.t226 VDD.t225 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X86 a_20090_158# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t48 VDD.t47 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X87 VSS.t40 a_30598_38# a_30498_n387# VSS.t39 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X88 a_1370_158# DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t301 VDD.t300 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X89 VSS.t232 PHI_1.t5 a_23030_n402# VSS.t231 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X90 a_26478_158# a_25962_n384# a_26330_n387# VSS.t49 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X91 a_35978_n384# a_35510_n402# VDD.t76 VDD.t75 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X92 a_36838_38# a_36494_158# VSS.t37 VSS.t36 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X93 a_n702_n387# a_n1930_n402# a_n946_158# VSS.t29 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X94 VDD.t162 a_30254_158# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t161 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X95 VDD.t102 a_36838_38# a_36698_158# VDD.t101 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X96 VDD.t6 a_58022_38# a_57882_158# VDD.t5 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X97 a_59143_n425# Q[10].t2 VSS.t286 VSS.t285 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X98 a_19722_n384# a_19254_n402# VDD.t72 VDD.t71 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X99 VSS.t85 a_24014_158# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t84 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X100 a_1002_n384# a_534_n402# VSS.t67 VSS.t66 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X101 gc[1].t0 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t110 VSS.t109 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X102 VDD.t145 PHI_1.t6 a_29270_n402# VDD.t144 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X103 a_39302_38# a_38958_158# VSS.t98 VSS.t97 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X104 VSS.t174 a_7758_158# Q[2].t0 VSS.t173 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X105 gc[5].t1 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t192 VDD.t191 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X106 a_36738_n387# a_35510_n402# a_36494_158# VSS.t76 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X107 a_8002_n387# a_6774_n402# a_7758_158# VSS.t202 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X108 a_17626_n387# Q[3].t2 VSS.t121 VSS.t120 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X109 a_33062_38# a_32718_158# VDD.t271 VDD.t270 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X110 a_36494_158# a_35510_n402# a_36346_158# VDD.t74 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X111 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[6].t3 VDD.t322 VDD.t321 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X112 a_30106_158# Q[5].t2 VDD.t324 VDD.t323 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X113 a_55066_n387# Q[9].t2 VSS.t323 VSS.t322 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X114 VDD.t337 a_11534_158# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t336 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X115 a_13850_158# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t78 VDD.t77 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X116 VDD.t172 a_39302_38# a_39162_158# VDD.t171 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X117 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t5 a_40423_n425# VSS.t235 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X118 a_14342_38# a_13998_158# VSS.t135 VSS.t134 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X119 a_18118_38# a_17774_158# VSS.t164 VSS.t163 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X120 VDD.t263 EN.t6 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t262 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X121 a_45442_n387# a_44214_n402# a_45198_158# VSS.t24 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X122 a_26330_n387# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t160 VSS.t159 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X123 VDD.t147 PHI_1.t7 a_54230_n402# VDD.t146 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X124 a_5638_38# a_5294_158# VDD.t19 VDD.t18 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X125 VDD.t125 a_45198_158# Q[8].t1 VDD.t124 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X126 a_14342_38# a_13998_158# VDD.t133 VDD.t132 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X127 a_13482_n384# a_13014_n402# VSS.t57 VSS.t56 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X128 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t7 a_59143_n425# VSS.t252 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X129 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[3].t3 VDD.t119 VDD.t118 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X130 a_18018_n387# a_16790_n402# a_17774_158# VSS.t310 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X131 a_24014_158# a_23030_n402# a_23866_158# VDD.t290 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X132 a_n742_158# a_n1462_n384# a_n946_158# VDD.t58 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X133 a_1518_158# a_1002_n384# a_1370_n387# VSS.t94 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X134 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t8 a_2983_n425# VSS.t253 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X135 a_5294_158# a_4778_n384# a_5146_n387# VSS.t79 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X136 a_30254_158# a_29270_n402# a_30106_158# VDD.t280 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X137 gc[4].t0 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t278 VSS.t277 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X138 VSS.t168 a_39302_38# a_39202_n387# VSS.t167 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X139 gc[9].t1 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t121 VDD.t120 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X140 a_15463_n425# Q[3].t4 VSS.t268 VSS.t267 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X141 gc[3].t0 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t312 VSS.t311 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X142 VSS.t137 a_26478_158# Q[5].t0 VSS.t136 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X143 a_30598_38# a_30254_158# VSS.t156 VSS.t155 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X144 VDD.t112 PHI_2.t6 a_534_n402# VDD.t111 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X145 VSS.t143 PHI_1.t8 a_4310_n402# VSS.t142 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X146 VDD.t182 PHI_1.t9 a_35510_n402# VDD.t181 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X147 a_36838_38# a_36494_158# VDD.t37 VDD.t36 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X148 a_45402_158# a_44682_n384# a_45198_158# VDD.t287 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X149 a_57530_158# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t69 VDD.t68 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X150 a_4778_n384# a_4310_n402# VSS.t152 VSS.t151 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X151 VDD.t135 a_26478_158# Q[5].t1 VDD.t134 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X152 a_52903_n425# Q[9].t3 VSS.t2 VSS.t1 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X153 a_n946_158# a_n1930_n402# a_n1094_158# VDD.t29 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X154 a_36698_158# a_35978_n384# a_36494_158# VDD.t73 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X155 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[7].t3 VDD.t194 VDD.t193 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X156 a_7610_158# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t286 VDD.t285 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X157 a_13998_158# a_13014_n402# a_13850_158# VDD.t55 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X158 a_38958_158# a_38442_n384# a_38810_n387# VSS.t321 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X159 a_45198_158# a_44682_n384# a_45050_n387# VSS.t281 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X160 VDD.t114 PHI_2.t7 a_6774_n402# VDD.t113 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X161 VSS.t204 PHI_2.t8 a_6774_n402# VSS.t203 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X162 a_48458_n384# a_47990_n402# VDD.t11 VDD.t10 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X163 gc[6].t1 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t307 VDD.t306 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X164 a_58022_38# a_57678_158# VSS.t189 VSS.t188 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X165 VSS.t199 a_51782_38# a_51682_n387# VSS.t198 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X166 VDD.t309 a_5638_38# a_5498_158# VDD.t308 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X167 a_18118_38# a_17774_158# VDD.t168 VDD.t167 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X168 VDD.t176 a_51438_158# Q[9].t1 VDD.t175 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X169 VSS.t206 PHI_2.t9 a_44214_n402# VSS.t205 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X170 a_55458_n387# a_54230_n402# a_55214_158# VSS.t192 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X171 a_n1094_158# D_in.t1 VDD.t210 VDD.t209 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X172 a_17774_158# a_17258_n384# a_17626_n387# VSS.t264 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X173 a_20238_158# a_19722_n384# a_20090_n387# VSS.t313 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X174 a_36346_n387# Q[6].t4 VSS.t316 VSS.t315 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X175 VDD.t208 a_45542_38# a_45402_158# VDD.t207 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X176 a_7610_n387# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t280 VSS.t279 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X177 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t9 a_15463_n425# VSS.t246 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X178 VDD.t257 EN.t10 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t256 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X179 a_30458_158# a_29738_n384# a_30254_158# VDD.t117 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X180 a_42586_158# Q[7].t4 VDD.t196 VDD.t195 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X181 a_50922_n384# a_50454_n402# VDD.t46 VDD.t45 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X182 a_1862_38# a_1518_158# VDD.t15 VDD.t14 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X183 VDD.t184 PHI_1.t10 a_16790_n402# VDD.t183 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X184 a_23498_n384# a_23030_n402# VSS.t283 VSS.t282 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X185 VDD.t217 PHI_2.t10 a_37974_n402# VDD.t216 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X186 a_57678_158# a_56694_n402# a_57530_158# VDD.t218 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X187 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t11 a_52903_n425# VSS.t247 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X188 a_14202_158# a_13482_n384# a_13998_158# VDD.t318 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X189 gc[3].t1 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t316 VDD.t315 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X190 VSS.t178 PHI_1.t11 a_16790_n402# VSS.t177 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X191 a_26330_158# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t164 VDD.t163 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X192 a_33062_38# a_32718_158# VSS.t261 VSS.t260 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X193 a_57922_n387# a_56694_n402# a_57678_158# VSS.t213 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X194 VSS.t19 a_5294_158# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t18 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X195 a_20582_38# a_20238_158# VDD.t60 VDD.t59 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X196 gc[10].t0 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t51 VSS.t50 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X197 VDD.t230 a_8102_38# a_7962_158# VDD.t229 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X198 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[4].t4 VDD.t248 VDD.t247 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X199 a_42218_n384# a_41750_n402# VDD.t129 VDD.t128 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X200 a_1762_n387# a_534_n402# a_1518_158# VSS.t65 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X201 a_7758_158# a_6774_n402# a_7610_158# VDD.t213 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X202 a_25962_n384# a_25494_n402# VDD.t154 VDD.t153 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X203 VSS.t106 a_49318_38# a_49218_n387# VSS.t105 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X204 VDD.t139 a_26822_38# a_26682_158# VDD.t138 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X205 VSS.t251 PHI_2.t11 a_25494_n402# VSS.t250 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X206 a_25962_n384# a_25494_n402# VSS.t149 VSS.t148 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X207 a_32202_n384# a_31734_n402# VSS.t43 VSS.t42 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X208 a_11878_38# a_11534_158# VSS.t329 VSS.t328 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X209 a_17258_n384# a_16790_n402# VDD.t314 VDD.t313 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X210 VDD.t240 PHI_1.t12 a_41750_n402# VDD.t239 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X211 a_43078_38# a_42734_158# VDD.t305 VDD.t304 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X212 VDD.t259 PHI_2.t12 a_19254_n402# VDD.t258 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X213 VDD.t269 a_32718_158# Q[6].t1 VDD.t268 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X214 gc[6].t0 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t303 VSS.t302 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X215 VSS.t4 a_58022_38# a_57922_n387# VSS.t3 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X216 VDD.t93 a_n602_38# a_n742_158# VDD.t92 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X217 a_27943_n425# Q[5].t3 VSS.t318 VSS.t317 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X218 a_34183_n425# Q[6].t5 VSS.t276 VSS.t275 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X219 VSS.t96 a_38958_158# Q[7].t0 VSS.t95 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X220 VSS.t127 a_45198_158# Q[8].t0 VSS.t126 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X221 VDD.t279 a_18118_38# a_17978_158# VDD.t278 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X222 a_55214_158# a_54698_n384# a_55066_n387# VSS.t0 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X223 a_57882_158# a_57162_n384# a_57678_158# VDD.t158 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X224 a_51438_158# a_50454_n402# a_51290_158# VDD.t44 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X225 a_20090_n387# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t48 VSS.t47 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X226 a_11778_n387# a_10550_n402# a_11534_158# VSS.t195 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X227 VDD.t242 PHI_1.t13 a_4310_n402# VDD.t241 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X228 gc[7].t1 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t87 VDD.t86 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X229 a_57678_158# a_57162_n384# a_57530_n387# VSS.t154 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X230 a_58022_38# a_57678_158# VDD.t200 VDD.t199 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X231 VDD.t149 a_55214_158# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t148 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X232 a_49178_158# a_48458_n384# a_48974_158# VDD.t293 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X233 a_7962_158# a_7242_n384# a_7758_158# VDD.t126 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X234 a_11386_158# Q[2].t2 VDD.t143 VDD.t142 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X235 VDD.t261 PHI_2.t13 a_44214_n402# VDD.t260 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X236 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[10].t3 VDD.t292 VDD.t291 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X237 VSS.t237 PHI_1.t14 a_54230_n402# VSS.t236 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X238 a_1518_158# a_534_n402# a_1370_158# VDD.t65 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X239 VSS.t162 a_17774_158# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t161 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X240 VSS.t60 a_20238_158# Q[4].t0 VSS.t59 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X241 a_24358_38# a_24014_158# VDD.t85 VDD.t84 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X242 a_26478_158# a_25494_n402# a_26330_158# VDD.t152 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X243 VSS.t81 a_33062_38# a_32962_n387# VSS.t80 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X244 VDD.t131 a_13998_158# Q[3].t1 VDD.t130 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X245 a_5638_38# a_5294_158# VSS.t17 VSS.t16 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X246 a_20482_n387# a_19254_n402# a_20238_158# VSS.t72 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X247 VDD.t212 a_51782_38# a_51642_158# VDD.t211 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X248 a_n602_38# a_n946_158# VSS.t33 VSS.t32 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X249 gc[1].t1 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t104 VDD.t103 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X250 VDD.t186 EN.t12 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t185 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X251 a_36494_158# a_35978_n384# a_36346_n387# VSS.t73 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X252 a_32718_158# a_32202_n384# a_32570_n387# VSS.t258 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X253 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t13 a_34183_n425# VSS.t179 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X254 a_48826_n387# Q[8].t2 VSS.t293 VSS.t292 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X255 a_51642_158# a_50922_n384# a_51438_158# VDD.t277 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X256 VDD.t35 a_36494_158# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t34 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X257 a_39302_38# a_38958_158# VDD.t98 VDD.t97 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X258 a_n1462_n384# a_n1930_n402# VDD.t28 VDD.t27 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X259 VDD.t326 PHI_2.t14 a_25494_n402# VDD.t325 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X260 VDD.t21 a_43078_38# a_42938_158# VDD.t20 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X261 a_48826_158# Q[8].t3 VDD.t297 VDD.t296 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X262 VSS.t100 PHI_1.t15 a_35510_n402# VSS.t99 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X263 a_35978_n384# a_35510_n402# VSS.t75 VSS.t74 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X264 a_42218_n384# a_41750_n402# VSS.t131 VSS.t130 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X265 a_49318_38# a_48974_158# VSS.t223 VSS.t222 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X266 a_1722_158# a_1002_n384# a_1518_158# VDD.t94 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X267 VSS.t26 a_14342_38# a_14242_n387# VSS.t25 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X268 a_26682_158# a_25962_n384# a_26478_158# VDD.t49 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X269 a_57530_n387# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t69 VSS.t68 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X270 a_51782_38# a_51438_158# VSS.t172 VSS.t171 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X271 a_45542_38# a_45198_158# VSS.t125 VSS.t124 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X272 a_20238_158# a_19254_n402# a_20090_158# VDD.t70 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X273 a_11534_158# a_11018_n384# a_11386_n387# VSS.t259 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X274 a_54698_n384# a_54230_n402# VDD.t202 VDD.t201 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X275 a_5146_158# Q[1].t4 VDD.t190 VDD.t189 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X276 a_1370_n387# DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t297 VSS.t296 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X277 VDD.t188 EN.t14 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t187 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X278 a_38442_n384# a_37974_n402# VDD.t53 VDD.t52 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X279 a_44682_n384# a_44214_n402# VSS.t23 VSS.t22 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X280 a_n602_38# a_n946_158# VDD.t31 VDD.t30 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X281 VDD.t166 a_17774_158# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t165 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X282 VSS.t102 PHI_1.t16 a_n1930_n402# VSS.t101 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X283 a_4778_n384# a_4310_n402# VDD.t157 VDD.t156 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X284 VSS.t305 a_5638_38# a_5538_n387# VSS.t304 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X285 VSS.t104 PHI_1.t17 a_10550_n402# VSS.t103 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X286 a_13998_158# a_13482_n384# a_13850_n387# VSS.t314 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X287 VDD.t89 a_24358_38# a_24218_158# VDD.t88 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X288 a_24358_38# a_24014_158# VSS.t83 VSS.t82 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X289 a_30598_38# a_30254_158# VDD.t160 VDD.t159 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X290 a_30106_n387# Q[5].t4 VSS.t91 VSS.t90 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X291 a_48974_158# a_47990_n402# a_48826_158# VDD.t9 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X292 gc[9].t0 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t123 VSS.t122 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X293 VSS.t187 a_57678_158# Q[10].t0 VSS.t186 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X294 gc[10].t1 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t51 VDD.t50 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X295 a_46663_n425# Q[8].t4 VSS.t295 VSS.t294 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X296 VSS.t21 a_43078_38# a_42978_n387# VSS.t20 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X297 VDD.t13 a_1518_158# Q[1].t1 VDD.t12 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X298 VSS.t11 a_1518_158# Q[1].t0 VSS.t10 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X299 VDD.t244 EN.t15 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t243 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X300 a_38810_n387# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t291 VSS.t290 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X301 VDD.t328 PHI_2.t15 a_50454_n402# VDD.t327 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X302 VSS.t31 a_n946_158# DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t30 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X303 a_20442_158# a_19722_n384# a_20238_158# VDD.t317 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X304 a_32570_158# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t170 VDD.t169 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X305 a_30498_n387# a_29270_n402# a_30254_158# VSS.t272 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X306 a_5294_158# a_4310_n402# a_5146_158# VDD.t155 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X307 a_7242_n384# a_6774_n402# VSS.t201 VSS.t200 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X308 a_11386_n387# Q[2].t3 VSS.t255 VSS.t254 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X309 VDD.t303 a_42734_158# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t302 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X310 a_17626_158# Q[3].t5 VDD.t276 VDD.t275 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X311 VSS.t35 a_36494_158# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t34 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X312 VSS.t93 a_n602_38# a_n702_n387# VSS.t92 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X313 a_32202_n384# a_31734_n402# VDD.t42 VDD.t41 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X314 a_n1462_n384# a_n1930_n402# VSS.t28 VSS.t27 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X315 a_32962_n387# a_31734_n402# a_32718_158# VSS.t41 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X316 a_9223_n425# Q[2].t4 VSS.t257 VSS.t256 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X317 a_13850_n387# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t78 VSS.t77 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X318 a_23498_n384# a_23030_n402# VDD.t289 VDD.t288 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X319 a_42734_158# a_41750_n402# a_42586_158# VDD.t127 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X320 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[8].t5 VDD.t299 VDD.t298 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X321 a_45542_38# a_45198_158# VDD.t123 VDD.t122 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X322 VDD.t330 PHI_2.t16 a_31734_n402# VDD.t329 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X323 a_48974_158# a_48458_n384# a_48826_n387# VSS.t287 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X324 VSS.t89 a_24358_38# a_24258_n387# VSS.t88 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X325 a_51438_158# a_50922_n384# a_51290_n387# VSS.t269 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X326 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t16 a_46663_n425# VSS.t238 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X327 VSS.t327 a_11534_158# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t326 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X328 a_17258_n384# a_16790_n402# VSS.t309 VSS.t308 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X329 VDD.t246 EN.t17 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t245 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X330 a_17774_158# a_16790_n402# a_17626_158# VDD.t312 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X331 a_54698_n384# a_54230_n402# VSS.t191 VSS.t190 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X332 VDD.t17 a_5294_158# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t16 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X333 a_8102_38# a_7758_158# VDD.t178 VDD.t177 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X334 VDD.t232 EN.t18 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t231 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X335 VSS.t141 a_26822_38# a_26722_n387# VSS.t140 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X336 VDD.t198 a_57678_158# Q[10].t1 VDD.t197 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X337 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[2].t5 VDD.t265 VDD.t264 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X338 VSS.t133 a_13998_158# Q[3].t0 VSS.t132 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X339 VDD.t253 PHI_1.t18 a_23030_n402# VDD.t252 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X340 a_39162_158# a_38442_n384# a_38958_158# VDD.t333 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X341 a_11018_n384# a_10550_n402# VDD.t206 VDD.t205 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X342 VSS.t208 PHI_2.t17 a_19254_n402# VSS.t207 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X343 a_19722_n384# a_19254_n402# VSS.t71 VSS.t70 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X344 VDD.t83 a_24014_158# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t82 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X345 a_24014_158# a_23498_n384# a_23866_n387# VSS.t38 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X346 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[5].t5 VDD.t91 VDD.t90 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X347 a_30254_158# a_29738_n384# a_30106_n387# VSS.t119 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X348 VDD.t40 a_30598_38# a_30458_158# VDD.t39 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X349 VSS.t210 PHI_2.t18 a_56694_n402# VSS.t209 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X350 VDD.t335 a_1862_38# a_1722_158# VDD.t334 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X351 a_5498_158# a_4778_n384# a_5294_158# VDD.t79 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X352 a_43078_38# a_42734_158# VSS.t299 VSS.t298 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X353 gc[4].t1 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t284 VDD.t283 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X354 a_39202_n387# a_37974_n402# a_38958_158# VSS.t52 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X355 a_49318_38# a_48974_158# VDD.t222 VDD.t221 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X356 a_11534_158# a_10550_n402# a_11386_158# VDD.t204 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X357 VDD.t96 a_38958_158# Q[7].t1 VDD.t95 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X358 a_42938_158# a_42218_n384# a_42734_158# VDD.t249 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X359 a_55066_158# Q[9].t4 VDD.t4 VDD.t3 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X360 VSS.t212 PHI_2.t19 a_31734_n402# VSS.t211 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X361 a_2983_n425# Q[1].t5 VSS.t181 VSS.t180 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X362 VDD.t8 a_11878_38# a_11738_158# VDD.t7 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X363 VDD.t81 a_33062_38# a_32922_158# VDD.t80 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X364 a_38810_158# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t295 VDD.t294 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X365 a_42978_n387# a_41750_n402# a_42734_158# VSS.t129 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X366 VDD.t234 EN.t19 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t233 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X367 a_23866_n387# Q[4].t5 VSS.t15 VSS.t14 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X368 VDD.t255 PHI_1.t19 a_n1930_n402# VDD.t254 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X369 a_17978_158# a_17258_n384# a_17774_158# VDD.t272 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X370 a_14242_n387# a_13014_n402# a_13998_158# VSS.t55 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X371 VSS.t145 a_55214_158# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t144 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X372 VSS.t221 a_48974_158# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t220 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X373 a_40423_n425# Q[7].t5 VSS.t249 VSS.t248 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X374 a_44682_n384# a_44214_n402# VDD.t23 VDD.t22 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X375 VSS.t170 a_51438_158# Q[9].t0 VSS.t169 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X376 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[9].t5 VDD.t2 VDD.t1 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X377 a_51782_38# a_51438_158# VDD.t174 VDD.t173 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X378 a_11018_n384# a_10550_n402# VSS.t194 VSS.t193 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X379 a_51682_n387# a_50454_n402# a_51438_158# VSS.t44 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
R0 VSS.n59 VSS.t50 2230.39
R1 VSS.n52 VSS.t122 2226.52
R2 VSS.n45 VSS.t306 2226.52
R3 VSS.n38 VSS.t86 2226.52
R4 VSS.n31 VSS.t302 2226.52
R5 VSS.n24 VSS.t182 2226.52
R6 VSS.n17 VSS.t277 2226.52
R7 VSS.n10 VSS.t311 2226.52
R8 VSS.n3 VSS.t111 2226.52
R9 VSS.t109 VSS.n178 2226.52
R10 VSS.t186 VSS.t188 2202.58
R11 VSS.t68 VSS.t214 2202.58
R12 VSS.t144 VSS.t146 2202.58
R13 VSS.t322 VSS.t190 2202.58
R14 VSS.t169 VSS.t171 2202.58
R15 VSS.t63 VSS.t45 2202.58
R16 VSS.t220 VSS.t222 2202.58
R17 VSS.t292 VSS.t7 2202.58
R18 VSS.t126 VSS.t124 2202.58
R19 VSS.t265 VSS.t22 2202.58
R20 VSS.t300 VSS.t298 2202.58
R21 VSS.t184 VSS.t130 2202.58
R22 VSS.t95 VSS.t97 2202.58
R23 VSS.t290 VSS.t53 2202.58
R24 VSS.t34 VSS.t36 2202.58
R25 VSS.t315 VSS.t74 2202.58
R26 VSS.t262 VSS.t260 2202.58
R27 VSS.t165 VSS.t42 2202.58
R28 VSS.t157 VSS.t155 2202.58
R29 VSS.t90 VSS.t273 2202.58
R30 VSS.t136 VSS.t138 2202.58
R31 VSS.t159 VSS.t148 2202.58
R32 VSS.t84 VSS.t82 2202.58
R33 VSS.t14 VSS.t282 2202.58
R34 VSS.t59 VSS.t61 2202.58
R35 VSS.t47 VSS.t70 2202.58
R36 VSS.t161 VSS.t163 2202.58
R37 VSS.t120 VSS.t308 2202.58
R38 VSS.t132 VSS.t134 2202.58
R39 VSS.t77 VSS.t56 2202.58
R40 VSS.t326 VSS.t328 2202.58
R41 VSS.t254 VSS.t193 2202.58
R42 VSS.t173 VSS.t175 2202.58
R43 VSS.t279 VSS.t200 2202.58
R44 VSS.t16 VSS.t18 2202.58
R45 VSS.t151 VSS.t227 2202.58
R46 VSS.t12 VSS.t10 2202.58
R47 VSS.t66 VSS.t296 2202.58
R48 VSS.t32 VSS.t30 2202.58
R49 VSS.t27 VSS.t288 2202.58
R50 VSS.n53 VSS.n52 1819.52
R51 VSS.n46 VSS.n45 1819.52
R52 VSS.n39 VSS.n38 1819.52
R53 VSS.n32 VSS.n31 1819.52
R54 VSS.n25 VSS.n24 1819.52
R55 VSS.n18 VSS.n17 1819.52
R56 VSS.n11 VSS.n10 1819.52
R57 VSS.n4 VSS.n3 1819.52
R58 VSS.n178 VSS.n177 1819.52
R59 VSS.n56 VSS.t144 1747.7
R60 VSS.n49 VSS.t220 1747.7
R61 VSS.n42 VSS.t300 1747.7
R62 VSS.n35 VSS.t34 1747.7
R63 VSS.n28 VSS.t157 1747.7
R64 VSS.n21 VSS.t84 1747.7
R65 VSS.n14 VSS.t161 1747.7
R66 VSS.n7 VSS.t326 1747.7
R67 VSS.t18 VSS.n176 1747.7
R68 VSS.t30 VSS.n181 1747.7
R69 VSS.t3 VSS.t213 1556.17
R70 VSS.t214 VSS.t209 1556.17
R71 VSS.t319 VSS.t192 1556.17
R72 VSS.t190 VSS.t236 1556.17
R73 VSS.t198 VSS.t44 1556.17
R74 VSS.t45 VSS.t117 1556.17
R75 VSS.t105 VSS.t9 1556.17
R76 VSS.t7 VSS.t229 1556.17
R77 VSS.t196 VSS.t24 1556.17
R78 VSS.t22 VSS.t205 1556.17
R79 VSS.t20 VSS.t129 1556.17
R80 VSS.t130 VSS.t244 1556.17
R81 VSS.t167 VSS.t52 1556.17
R82 VSS.t53 VSS.t218 1556.17
R83 VSS.t107 VSS.t76 1556.17
R84 VSS.t74 VSS.t99 1556.17
R85 VSS.t80 VSS.t41 1556.17
R86 VSS.t42 VSS.t211 1556.17
R87 VSS.t39 VSS.t272 1556.17
R88 VSS.t273 VSS.t242 1556.17
R89 VSS.t140 VSS.t150 1556.17
R90 VSS.t148 VSS.t250 1556.17
R91 VSS.t88 VSS.t284 1556.17
R92 VSS.t282 VSS.t231 1556.17
R93 VSS.t113 VSS.t72 1556.17
R94 VSS.t70 VSS.t207 1556.17
R95 VSS.t270 VSS.t310 1556.17
R96 VSS.t308 VSS.t177 1556.17
R97 VSS.t25 VSS.t55 1556.17
R98 VSS.t56 VSS.t115 1556.17
R99 VSS.t5 VSS.t195 1556.17
R100 VSS.t193 VSS.t103 1556.17
R101 VSS.t233 VSS.t202 1556.17
R102 VSS.t200 VSS.t203 1556.17
R103 VSS.t153 VSS.t304 1556.17
R104 VSS.t142 VSS.t151 1556.17
R105 VSS.t65 VSS.t324 1556.17
R106 VSS.t216 VSS.t66 1556.17
R107 VSS.t29 VSS.t92 1556.17
R108 VSS.t101 VSS.t27 1556.17
R109 VSS VSS.t252 1550.18
R110 VSS VSS.t247 1550.18
R111 VSS VSS.t238 1550.18
R112 VSS VSS.t235 1550.18
R113 VSS VSS.t179 1550.18
R114 VSS VSS.t224 1550.18
R115 VSS VSS.t225 1550.18
R116 VSS VSS.t246 1550.18
R117 VSS VSS.t226 1550.18
R118 VSS.t253 VSS 1550.18
R119 VSS VSS.t186 1508.29
R120 VSS VSS.t169 1508.29
R121 VSS VSS.t126 1508.29
R122 VSS VSS.t95 1508.29
R123 VSS VSS.t262 1508.29
R124 VSS VSS.t136 1508.29
R125 VSS VSS.t59 1508.29
R126 VSS VSS.t132 1508.29
R127 VSS VSS.t173 1508.29
R128 VSS.t10 VSS 1508.29
R129 VSS.t188 VSS.t3 1340.7
R130 VSS.t213 VSS.t154 1340.7
R131 VSS.t146 VSS.t319 1340.7
R132 VSS.t192 VSS.t0 1340.7
R133 VSS.t171 VSS.t198 1340.7
R134 VSS.t44 VSS.t269 1340.7
R135 VSS.t222 VSS.t105 1340.7
R136 VSS.t9 VSS.t287 1340.7
R137 VSS.t124 VSS.t196 1340.7
R138 VSS.t24 VSS.t281 1340.7
R139 VSS.t298 VSS.t20 1340.7
R140 VSS.t129 VSS.t241 1340.7
R141 VSS.t97 VSS.t167 1340.7
R142 VSS.t52 VSS.t321 1340.7
R143 VSS.t36 VSS.t107 1340.7
R144 VSS.t76 VSS.t73 1340.7
R145 VSS.t260 VSS.t80 1340.7
R146 VSS.t41 VSS.t258 1340.7
R147 VSS.t155 VSS.t39 1340.7
R148 VSS.t272 VSS.t119 1340.7
R149 VSS.t138 VSS.t140 1340.7
R150 VSS.t150 VSS.t49 1340.7
R151 VSS.t82 VSS.t88 1340.7
R152 VSS.t284 VSS.t38 1340.7
R153 VSS.t61 VSS.t113 1340.7
R154 VSS.t72 VSS.t313 1340.7
R155 VSS.t163 VSS.t270 1340.7
R156 VSS.t310 VSS.t264 1340.7
R157 VSS.t134 VSS.t25 1340.7
R158 VSS.t55 VSS.t314 1340.7
R159 VSS.t328 VSS.t5 1340.7
R160 VSS.t195 VSS.t259 1340.7
R161 VSS.t175 VSS.t233 1340.7
R162 VSS.t202 VSS.t128 1340.7
R163 VSS.t304 VSS.t16 1340.7
R164 VSS.t79 VSS.t153 1340.7
R165 VSS.t324 VSS.t12 1340.7
R166 VSS.t94 VSS.t65 1340.7
R167 VSS.t92 VSS.t32 1340.7
R168 VSS.t58 VSS.t29 1340.7
R169 VSS.n184 VSS 1104.92
R170 VSS.t252 VSS.t285 1101.29
R171 VSS VSS.n56 1101.29
R172 VSS VSS.n53 1101.29
R173 VSS.t247 VSS.t1 1101.29
R174 VSS VSS.n49 1101.29
R175 VSS VSS.n46 1101.29
R176 VSS.t238 VSS.t294 1101.29
R177 VSS VSS.n42 1101.29
R178 VSS VSS.n39 1101.29
R179 VSS.t235 VSS.t248 1101.29
R180 VSS VSS.n35 1101.29
R181 VSS VSS.n32 1101.29
R182 VSS.t179 VSS.t275 1101.29
R183 VSS VSS.n28 1101.29
R184 VSS VSS.n25 1101.29
R185 VSS.t224 VSS.t317 1101.29
R186 VSS VSS.n21 1101.29
R187 VSS VSS.n18 1101.29
R188 VSS.t225 VSS.t239 1101.29
R189 VSS VSS.n14 1101.29
R190 VSS VSS.n11 1101.29
R191 VSS.t246 VSS.t267 1101.29
R192 VSS VSS.n7 1101.29
R193 VSS VSS.n4 1101.29
R194 VSS.t226 VSS.t256 1101.29
R195 VSS.n176 VSS 1101.29
R196 VSS.n177 VSS 1101.29
R197 VSS.t180 VSS.t253 1101.29
R198 VSS.n181 VSS 1101.29
R199 VSS.t154 VSS.t68 1005.52
R200 VSS.t0 VSS.t322 1005.52
R201 VSS.t269 VSS.t63 1005.52
R202 VSS.t287 VSS.t292 1005.52
R203 VSS.t281 VSS.t265 1005.52
R204 VSS.t241 VSS.t184 1005.52
R205 VSS.t321 VSS.t290 1005.52
R206 VSS.t73 VSS.t315 1005.52
R207 VSS.t258 VSS.t165 1005.52
R208 VSS.t119 VSS.t90 1005.52
R209 VSS.t49 VSS.t159 1005.52
R210 VSS.t38 VSS.t14 1005.52
R211 VSS.t313 VSS.t47 1005.52
R212 VSS.t264 VSS.t120 1005.52
R213 VSS.t314 VSS.t77 1005.52
R214 VSS.t259 VSS.t254 1005.52
R215 VSS.t128 VSS.t279 1005.52
R216 VSS.t227 VSS.t79 1005.52
R217 VSS.t296 VSS.t94 1005.52
R218 VSS.t288 VSS.t58 1005.52
R219 VSS.t285 VSS 700.277
R220 VSS.t1 VSS 700.277
R221 VSS.t294 VSS 700.277
R222 VSS.t248 VSS 700.277
R223 VSS.t275 VSS 700.277
R224 VSS.t317 VSS 700.277
R225 VSS.t239 VSS 700.277
R226 VSS.t267 VSS 700.277
R227 VSS.t256 VSS 700.277
R228 VSS VSS.t180 700.277
R229 VSS.t50 VSS 694.292
R230 VSS.t209 VSS 694.292
R231 VSS.t236 VSS 694.292
R232 VSS.t122 VSS 694.292
R233 VSS.t117 VSS 694.292
R234 VSS.t229 VSS 694.292
R235 VSS.t306 VSS 694.292
R236 VSS.t205 VSS 694.292
R237 VSS.t244 VSS 694.292
R238 VSS.t86 VSS 694.292
R239 VSS.t218 VSS 694.292
R240 VSS.t99 VSS 694.292
R241 VSS.t302 VSS 694.292
R242 VSS.t211 VSS 694.292
R243 VSS.t242 VSS 694.292
R244 VSS.t182 VSS 694.292
R245 VSS.t250 VSS 694.292
R246 VSS.t231 VSS 694.292
R247 VSS.t277 VSS 694.292
R248 VSS.t207 VSS 694.292
R249 VSS.t177 VSS 694.292
R250 VSS.t311 VSS 694.292
R251 VSS.t115 VSS 694.292
R252 VSS.t103 VSS 694.292
R253 VSS.t111 VSS 694.292
R254 VSS.t203 VSS 694.292
R255 VSS VSS.t142 694.292
R256 VSS VSS.t109 694.292
R257 VSS VSS.t216 694.292
R258 VSS VSS.t101 694.292
R259 VSS.n63 VSS.t69 8.79702
R260 VSS.n68 VSS.t323 8.79702
R261 VSS.n76 VSS.t64 8.79702
R262 VSS.n81 VSS.t293 8.79702
R263 VSS.n89 VSS.t266 8.79702
R264 VSS.n94 VSS.t185 8.79702
R265 VSS.n102 VSS.t291 8.79702
R266 VSS.n107 VSS.t316 8.79702
R267 VSS.n115 VSS.t166 8.79702
R268 VSS.n120 VSS.t91 8.79702
R269 VSS.n128 VSS.t160 8.79702
R270 VSS.n133 VSS.t15 8.79702
R271 VSS.n141 VSS.t48 8.79702
R272 VSS.n146 VSS.t121 8.79702
R273 VSS.n154 VSS.t78 8.79702
R274 VSS.n159 VSS.t255 8.79702
R275 VSS.n167 VSS.t280 8.79702
R276 VSS.n172 VSS.t228 8.79702
R277 VSS.n191 VSS.t297 8.79702
R278 VSS.n186 VSS.t289 8.79702
R279 VSS.n64 VSS.n57 6.40811
R280 VSS.n69 VSS.n54 6.40811
R281 VSS.n77 VSS.n50 6.40811
R282 VSS.n82 VSS.n47 6.40811
R283 VSS.n90 VSS.n43 6.40811
R284 VSS.n95 VSS.n40 6.40811
R285 VSS.n103 VSS.n36 6.40811
R286 VSS.n108 VSS.n33 6.40811
R287 VSS.n116 VSS.n29 6.40811
R288 VSS.n121 VSS.n26 6.40811
R289 VSS.n129 VSS.n22 6.40811
R290 VSS.n134 VSS.n19 6.40811
R291 VSS.n142 VSS.n15 6.40811
R292 VSS.n147 VSS.n12 6.40811
R293 VSS.n155 VSS.n8 6.40811
R294 VSS.n160 VSS.n5 6.40811
R295 VSS.n168 VSS.n1 6.40811
R296 VSS.n171 VSS.n170 6.40811
R297 VSS.n190 VSS.n180 6.40811
R298 VSS.n185 VSS.n183 6.40811
R299 VSS.n62 VSS.n58 6.4042
R300 VSS.n67 VSS.n55 6.4042
R301 VSS.n75 VSS.n51 6.4042
R302 VSS.n80 VSS.n48 6.4042
R303 VSS.n88 VSS.n44 6.4042
R304 VSS.n93 VSS.n41 6.4042
R305 VSS.n101 VSS.n37 6.4042
R306 VSS.n106 VSS.n34 6.4042
R307 VSS.n114 VSS.n30 6.4042
R308 VSS.n119 VSS.n27 6.4042
R309 VSS.n127 VSS.n23 6.4042
R310 VSS.n132 VSS.n20 6.4042
R311 VSS.n140 VSS.n16 6.4042
R312 VSS.n145 VSS.n13 6.4042
R313 VSS.n153 VSS.n9 6.4042
R314 VSS.n158 VSS.n6 6.4042
R315 VSS.n166 VSS.n2 6.4042
R316 VSS.n173 VSS.n169 6.4042
R317 VSS.n192 VSS.n179 6.4042
R318 VSS.n187 VSS.n182 6.4042
R319 VSS.n59 VSS.t51 4.63989
R320 VSS.n61 VSS.t187 4.63989
R321 VSS.n66 VSS.t145 4.63989
R322 VSS.n72 VSS.t123 4.63989
R323 VSS.n74 VSS.t170 4.63989
R324 VSS.n79 VSS.t221 4.63989
R325 VSS.n85 VSS.t307 4.63989
R326 VSS.n87 VSS.t127 4.63989
R327 VSS.n92 VSS.t301 4.63989
R328 VSS.n98 VSS.t87 4.63989
R329 VSS.n100 VSS.t96 4.63989
R330 VSS.n105 VSS.t35 4.63989
R331 VSS.n111 VSS.t303 4.63989
R332 VSS.n113 VSS.t263 4.63989
R333 VSS.n118 VSS.t158 4.63989
R334 VSS.n124 VSS.t183 4.63989
R335 VSS.n126 VSS.t137 4.63989
R336 VSS.n131 VSS.t85 4.63989
R337 VSS.n137 VSS.t278 4.63989
R338 VSS.n139 VSS.t60 4.63989
R339 VSS.n144 VSS.t162 4.63989
R340 VSS.n150 VSS.t312 4.63989
R341 VSS.n152 VSS.t133 4.63989
R342 VSS.n157 VSS.t327 4.63989
R343 VSS.n163 VSS.t112 4.63989
R344 VSS.n165 VSS.t174 4.63989
R345 VSS.n174 VSS.t19 4.63989
R346 VSS.n195 VSS.t110 4.63989
R347 VSS.n193 VSS.t11 4.63989
R348 VSS.n188 VSS.t31 4.63989
R349 VSS.n60 VSS.t286 4.51271
R350 VSS.n73 VSS.t2 4.51271
R351 VSS.n86 VSS.t295 4.51271
R352 VSS.n99 VSS.t249 4.51271
R353 VSS.n112 VSS.t276 4.51271
R354 VSS.n125 VSS.t318 4.51271
R355 VSS.n138 VSS.t240 4.51271
R356 VSS.n151 VSS.t268 4.51271
R357 VSS.n164 VSS.t257 4.51271
R358 VSS.n194 VSS.t181 4.51271
R359 VSS.n57 VSS.t215 3.9605
R360 VSS.n54 VSS.t191 3.9605
R361 VSS.n50 VSS.t46 3.9605
R362 VSS.n47 VSS.t8 3.9605
R363 VSS.n43 VSS.t23 3.9605
R364 VSS.n40 VSS.t131 3.9605
R365 VSS.n36 VSS.t54 3.9605
R366 VSS.n33 VSS.t75 3.9605
R367 VSS.n29 VSS.t43 3.9605
R368 VSS.n26 VSS.t274 3.9605
R369 VSS.n22 VSS.t149 3.9605
R370 VSS.n19 VSS.t283 3.9605
R371 VSS.n15 VSS.t71 3.9605
R372 VSS.n12 VSS.t309 3.9605
R373 VSS.n8 VSS.t57 3.9605
R374 VSS.n5 VSS.t194 3.9605
R375 VSS.n1 VSS.t201 3.9605
R376 VSS.n170 VSS.t152 3.9605
R377 VSS.n180 VSS.t67 3.9605
R378 VSS.n183 VSS.t28 3.9605
R379 VSS.n189 VSS.n181 3.6294
R380 VSS.n196 VSS.n178 3.6294
R381 VSS.n177 VSS.n0 3.6294
R382 VSS.n176 VSS.n175 3.6294
R383 VSS.n162 VSS.n3 3.6294
R384 VSS.n161 VSS.n4 3.6294
R385 VSS.n156 VSS.n7 3.6294
R386 VSS.n149 VSS.n10 3.6294
R387 VSS.n148 VSS.n11 3.6294
R388 VSS.n143 VSS.n14 3.6294
R389 VSS.n136 VSS.n17 3.6294
R390 VSS.n135 VSS.n18 3.6294
R391 VSS.n130 VSS.n21 3.6294
R392 VSS.n123 VSS.n24 3.6294
R393 VSS.n122 VSS.n25 3.6294
R394 VSS.n117 VSS.n28 3.6294
R395 VSS.n110 VSS.n31 3.6294
R396 VSS.n109 VSS.n32 3.6294
R397 VSS.n104 VSS.n35 3.6294
R398 VSS.n97 VSS.n38 3.6294
R399 VSS.n96 VSS.n39 3.6294
R400 VSS.n91 VSS.n42 3.6294
R401 VSS.n84 VSS.n45 3.6294
R402 VSS.n83 VSS.n46 3.6294
R403 VSS.n78 VSS.n49 3.6294
R404 VSS.n71 VSS.n52 3.6294
R405 VSS.n70 VSS.n53 3.6294
R406 VSS.n65 VSS.n56 3.6294
R407 VSS.n58 VSS.t189 2.07392
R408 VSS.n58 VSS.t4 2.07392
R409 VSS.n55 VSS.t147 2.07392
R410 VSS.n55 VSS.t320 2.07392
R411 VSS.n51 VSS.t172 2.07392
R412 VSS.n51 VSS.t199 2.07392
R413 VSS.n48 VSS.t223 2.07392
R414 VSS.n48 VSS.t106 2.07392
R415 VSS.n44 VSS.t125 2.07392
R416 VSS.n44 VSS.t197 2.07392
R417 VSS.n41 VSS.t299 2.07392
R418 VSS.n41 VSS.t21 2.07392
R419 VSS.n37 VSS.t98 2.07392
R420 VSS.n37 VSS.t168 2.07392
R421 VSS.n34 VSS.t37 2.07392
R422 VSS.n34 VSS.t108 2.07392
R423 VSS.n30 VSS.t261 2.07392
R424 VSS.n30 VSS.t81 2.07392
R425 VSS.n27 VSS.t156 2.07392
R426 VSS.n27 VSS.t40 2.07392
R427 VSS.n23 VSS.t139 2.07392
R428 VSS.n23 VSS.t141 2.07392
R429 VSS.n20 VSS.t83 2.07392
R430 VSS.n20 VSS.t89 2.07392
R431 VSS.n16 VSS.t62 2.07392
R432 VSS.n16 VSS.t114 2.07392
R433 VSS.n13 VSS.t164 2.07392
R434 VSS.n13 VSS.t271 2.07392
R435 VSS.n9 VSS.t135 2.07392
R436 VSS.n9 VSS.t26 2.07392
R437 VSS.n6 VSS.t329 2.07392
R438 VSS.n6 VSS.t6 2.07392
R439 VSS.n2 VSS.t176 2.07392
R440 VSS.n2 VSS.t234 2.07392
R441 VSS.n169 VSS.t17 2.07392
R442 VSS.n169 VSS.t305 2.07392
R443 VSS.n179 VSS.t13 2.07392
R444 VSS.n179 VSS.t325 2.07392
R445 VSS.n182 VSS.t33 2.07392
R446 VSS.n182 VSS.t93 2.07392
R447 VSS.n57 VSS.t210 1.84987
R448 VSS.n54 VSS.t237 1.84987
R449 VSS.n50 VSS.t118 1.84987
R450 VSS.n47 VSS.t230 1.84987
R451 VSS.n43 VSS.t206 1.84987
R452 VSS.n40 VSS.t245 1.84987
R453 VSS.n36 VSS.t219 1.84987
R454 VSS.n33 VSS.t100 1.84987
R455 VSS.n29 VSS.t212 1.84987
R456 VSS.n26 VSS.t243 1.84987
R457 VSS.n22 VSS.t251 1.84987
R458 VSS.n19 VSS.t232 1.84987
R459 VSS.n15 VSS.t208 1.84987
R460 VSS.n12 VSS.t178 1.84987
R461 VSS.n8 VSS.t116 1.84987
R462 VSS.n5 VSS.t104 1.84987
R463 VSS.n1 VSS.t204 1.84987
R464 VSS.n170 VSS.t143 1.84987
R465 VSS.n180 VSS.t217 1.84987
R466 VSS.n183 VSS.t102 1.84987
R467 VSS.n63 VSS.n62 0.4385
R468 VSS.n68 VSS.n67 0.4385
R469 VSS.n76 VSS.n75 0.4385
R470 VSS.n81 VSS.n80 0.4385
R471 VSS.n89 VSS.n88 0.4385
R472 VSS.n94 VSS.n93 0.4385
R473 VSS.n102 VSS.n101 0.4385
R474 VSS.n107 VSS.n106 0.4385
R475 VSS.n115 VSS.n114 0.4385
R476 VSS.n120 VSS.n119 0.4385
R477 VSS.n128 VSS.n127 0.4385
R478 VSS.n133 VSS.n132 0.4385
R479 VSS.n141 VSS.n140 0.4385
R480 VSS.n146 VSS.n145 0.4385
R481 VSS.n154 VSS.n153 0.4385
R482 VSS.n159 VSS.n158 0.4385
R483 VSS.n167 VSS.n166 0.4385
R484 VSS.n173 VSS.n172 0.4385
R485 VSS.n192 VSS.n191 0.4385
R486 VSS.n187 VSS.n186 0.4385
R487 VSS.n62 VSS.n61 0.2965
R488 VSS.n67 VSS.n66 0.2965
R489 VSS.n75 VSS.n74 0.2965
R490 VSS.n80 VSS.n79 0.2965
R491 VSS.n88 VSS.n87 0.2965
R492 VSS.n93 VSS.n92 0.2965
R493 VSS.n101 VSS.n100 0.2965
R494 VSS.n106 VSS.n105 0.2965
R495 VSS.n114 VSS.n113 0.2965
R496 VSS.n119 VSS.n118 0.2965
R497 VSS.n127 VSS.n126 0.2965
R498 VSS.n132 VSS.n131 0.2965
R499 VSS.n140 VSS.n139 0.2965
R500 VSS.n145 VSS.n144 0.2965
R501 VSS.n153 VSS.n152 0.2965
R502 VSS.n158 VSS.n157 0.2965
R503 VSS.n166 VSS.n165 0.2965
R504 VSS.n174 VSS.n173 0.2965
R505 VSS.n193 VSS.n192 0.2965
R506 VSS.n188 VSS.n187 0.2965
R507 VSS.n60 VSS.n59 0.28
R508 VSS.n73 VSS.n72 0.28
R509 VSS.n86 VSS.n85 0.28
R510 VSS.n99 VSS.n98 0.28
R511 VSS.n112 VSS.n111 0.28
R512 VSS.n125 VSS.n124 0.28
R513 VSS.n138 VSS.n137 0.28
R514 VSS.n151 VSS.n150 0.28
R515 VSS.n164 VSS.n163 0.28
R516 VSS.n195 VSS.n194 0.28
R517 VSS.n72 VSS.n71 0.2405
R518 VSS.n85 VSS.n84 0.2405
R519 VSS.n98 VSS.n97 0.2405
R520 VSS.n111 VSS.n110 0.2405
R521 VSS.n124 VSS.n123 0.2405
R522 VSS.n137 VSS.n136 0.2405
R523 VSS.n150 VSS.n149 0.2405
R524 VSS.n163 VSS.n162 0.2405
R525 VSS.n196 VSS.n195 0.2405
R526 VSS.n65 VSS.n64 0.2085
R527 VSS.n78 VSS.n77 0.2085
R528 VSS.n91 VSS.n90 0.2085
R529 VSS.n104 VSS.n103 0.2085
R530 VSS.n117 VSS.n116 0.2085
R531 VSS.n130 VSS.n129 0.2085
R532 VSS.n143 VSS.n142 0.2085
R533 VSS.n156 VSS.n155 0.2085
R534 VSS.n175 VSS.n168 0.2085
R535 VSS.n190 VSS.n189 0.2085
R536 VSS.n64 VSS.n63 0.2025
R537 VSS.n69 VSS.n68 0.2025
R538 VSS.n77 VSS.n76 0.2025
R539 VSS.n82 VSS.n81 0.2025
R540 VSS.n90 VSS.n89 0.2025
R541 VSS.n95 VSS.n94 0.2025
R542 VSS.n103 VSS.n102 0.2025
R543 VSS.n108 VSS.n107 0.2025
R544 VSS.n116 VSS.n115 0.2025
R545 VSS.n121 VSS.n120 0.2025
R546 VSS.n129 VSS.n128 0.2025
R547 VSS.n134 VSS.n133 0.2025
R548 VSS.n142 VSS.n141 0.2025
R549 VSS.n147 VSS.n146 0.2025
R550 VSS.n155 VSS.n154 0.2025
R551 VSS.n160 VSS.n159 0.2025
R552 VSS.n168 VSS.n167 0.2025
R553 VSS.n172 VSS.n171 0.2025
R554 VSS.n191 VSS.n190 0.2025
R555 VSS.n186 VSS.n185 0.2025
R556 VSS.n70 VSS 0.1645
R557 VSS.n83 VSS 0.1645
R558 VSS.n96 VSS 0.1645
R559 VSS.n109 VSS 0.1645
R560 VSS.n122 VSS 0.1645
R561 VSS.n135 VSS 0.1645
R562 VSS.n148 VSS 0.1645
R563 VSS.n161 VSS 0.1645
R564 VSS VSS.n0 0.1645
R565 VSS VSS.n184 0.1645
R566 VSS.n66 VSS.n65 0.0885
R567 VSS.n79 VSS.n78 0.0885
R568 VSS.n92 VSS.n91 0.0885
R569 VSS.n105 VSS.n104 0.0885
R570 VSS.n118 VSS.n117 0.0885
R571 VSS.n131 VSS.n130 0.0885
R572 VSS.n144 VSS.n143 0.0885
R573 VSS.n157 VSS.n156 0.0885
R574 VSS.n175 VSS.n174 0.0885
R575 VSS.n189 VSS.n188 0.0885
R576 VSS VSS.n70 0.0765
R577 VSS.n71 VSS 0.0765
R578 VSS VSS.n83 0.0765
R579 VSS.n84 VSS 0.0765
R580 VSS VSS.n96 0.0765
R581 VSS.n97 VSS 0.0765
R582 VSS VSS.n109 0.0765
R583 VSS.n110 VSS 0.0765
R584 VSS VSS.n122 0.0765
R585 VSS.n123 VSS 0.0765
R586 VSS VSS.n135 0.0765
R587 VSS.n136 VSS 0.0765
R588 VSS VSS.n148 0.0765
R589 VSS.n149 VSS 0.0765
R590 VSS VSS.n161 0.0765
R591 VSS.n162 VSS 0.0765
R592 VSS VSS.n0 0.0765
R593 VSS VSS.n196 0.0765
R594 VSS.n184 VSS 0.0765
R595 VSS.n61 VSS.n60 0.073
R596 VSS.n74 VSS.n73 0.073
R597 VSS.n87 VSS.n86 0.073
R598 VSS.n100 VSS.n99 0.073
R599 VSS.n113 VSS.n112 0.073
R600 VSS.n126 VSS.n125 0.073
R601 VSS.n139 VSS.n138 0.073
R602 VSS.n152 VSS.n151 0.073
R603 VSS.n165 VSS.n164 0.073
R604 VSS.n194 VSS.n193 0.073
R605 VSS VSS.n69 0.0445
R606 VSS VSS.n82 0.0445
R607 VSS VSS.n95 0.0445
R608 VSS VSS.n108 0.0445
R609 VSS VSS.n121 0.0445
R610 VSS VSS.n134 0.0445
R611 VSS VSS.n147 0.0445
R612 VSS VSS.n160 0.0445
R613 VSS.n171 VSS 0.0445
R614 VSS.n185 VSS 0.0445
R615 VDD.t197 VDD.t199 667.707
R616 VDD.t148 VDD.t150 667.707
R617 VDD.t175 VDD.t173 667.707
R618 VDD.t223 VDD.t221 667.707
R619 VDD.t124 VDD.t122 667.707
R620 VDD.t302 VDD.t304 667.707
R621 VDD.t95 VDD.t97 667.707
R622 VDD.t34 VDD.t36 667.707
R623 VDD.t268 VDD.t270 667.707
R624 VDD.t161 VDD.t159 667.707
R625 VDD.t134 VDD.t136 667.707
R626 VDD.t82 VDD.t84 667.707
R627 VDD.t61 VDD.t59 667.707
R628 VDD.t165 VDD.t167 667.707
R629 VDD.t130 VDD.t132 667.707
R630 VDD.t336 VDD.t338 667.707
R631 VDD.t179 VDD.t177 667.707
R632 VDD.t18 VDD.t16 667.707
R633 VDD.t14 VDD.t12 667.707
R634 VDD.t30 VDD.t32 667.707
R635 VDD.t68 VDD.t219 574.104
R636 VDD.t3 VDD.t201 574.104
R637 VDD.t63 VDD.t45 574.104
R638 VDD.t296 VDD.t10 574.104
R639 VDD.t273 VDD.t22 574.104
R640 VDD.t195 VDD.t128 574.104
R641 VDD.t294 VDD.t52 574.104
R642 VDD.t319 VDD.t75 574.104
R643 VDD.t169 VDD.t41 574.104
R644 VDD.t323 VDD.t281 574.104
R645 VDD.t163 VDD.t153 574.104
R646 VDD.t140 VDD.t288 574.104
R647 VDD.t47 VDD.t71 574.104
R648 VDD.t275 VDD.t313 574.104
R649 VDD.t77 VDD.t56 574.104
R650 VDD.t142 VDD.t205 574.104
R651 VDD.t285 VDD.t214 574.104
R652 VDD.t156 VDD.t189 574.104
R653 VDD.t66 VDD.t300 574.104
R654 VDD.t27 VDD.t209 574.104
R655 VDD.n59 VDD.t50 569.532
R656 VDD.n52 VDD.t120 564.744
R657 VDD.n45 VDD.t310 564.744
R658 VDD.n38 VDD.t86 564.744
R659 VDD.n31 VDD.t306 564.744
R660 VDD.n24 VDD.t191 564.744
R661 VDD.n17 VDD.t283 564.744
R662 VDD.n10 VDD.t315 564.744
R663 VDD.n3 VDD.t105 564.744
R664 VDD.t103 VDD.n187 564.744
R665 VDD.n53 VDD.n52 474.26
R666 VDD.n46 VDD.n45 474.26
R667 VDD.n39 VDD.n38 474.26
R668 VDD.n32 VDD.n31 474.26
R669 VDD.n25 VDD.n24 474.26
R670 VDD.n18 VDD.n17 474.26
R671 VDD.n11 VDD.n10 474.26
R672 VDD.n4 VDD.n3 474.26
R673 VDD.n187 VDD.n186 474.26
R674 VDD.n56 VDD.t148 471.139
R675 VDD.n49 VDD.t223 471.139
R676 VDD.n42 VDD.t302 471.139
R677 VDD.n35 VDD.t34 471.139
R678 VDD.n28 VDD.t161 471.139
R679 VDD.n21 VDD.t82 471.139
R680 VDD.n14 VDD.t165 471.139
R681 VDD.n7 VDD.t336 471.139
R682 VDD.t16 VDD.n185 471.139
R683 VDD.t32 VDD.n190 471.139
R684 VDD VDD.t197 410.296
R685 VDD VDD.t175 410.296
R686 VDD VDD.t124 410.296
R687 VDD VDD.t95 410.296
R688 VDD VDD.t268 410.296
R689 VDD VDD.t134 410.296
R690 VDD VDD.t61 410.296
R691 VDD VDD.t130 410.296
R692 VDD VDD.t179 410.296
R693 VDD.t12 VDD 410.296
R694 VDD.t219 VDD.t115 405.616
R695 VDD.t201 VDD.t146 405.616
R696 VDD.t45 VDD.t327 405.616
R697 VDD.t10 VDD.t227 405.616
R698 VDD.t22 VDD.t260 405.616
R699 VDD.t128 VDD.t239 405.616
R700 VDD.t52 VDD.t216 405.616
R701 VDD.t75 VDD.t181 405.616
R702 VDD.t41 VDD.t329 405.616
R703 VDD.t281 VDD.t144 405.616
R704 VDD.t153 VDD.t325 405.616
R705 VDD.t288 VDD.t252 405.616
R706 VDD.t71 VDD.t258 405.616
R707 VDD.t313 VDD.t183 405.616
R708 VDD.t56 VDD.t109 405.616
R709 VDD.t205 VDD.t250 405.616
R710 VDD.t214 VDD.t113 405.616
R711 VDD.t241 VDD.t156 405.616
R712 VDD.t111 VDD.t66 405.616
R713 VDD.t254 VDD.t27 405.616
R714 VDD VDD.t233 390.017
R715 VDD VDD.t262 390.017
R716 VDD VDD.t235 390.017
R717 VDD VDD.t243 390.017
R718 VDD VDD.t185 390.017
R719 VDD VDD.t256 390.017
R720 VDD VDD.t231 390.017
R721 VDD VDD.t187 390.017
R722 VDD VDD.t237 390.017
R723 VDD.t245 VDD 390.017
R724 VDD.t5 VDD.t158 374.416
R725 VDD.t331 VDD.t0 374.416
R726 VDD.t211 VDD.t277 374.416
R727 VDD.t99 VDD.t293 374.416
R728 VDD.t207 VDD.t287 374.416
R729 VDD.t20 VDD.t249 374.416
R730 VDD.t171 VDD.t333 374.416
R731 VDD.t101 VDD.t73 374.416
R732 VDD.t80 VDD.t266 374.416
R733 VDD.t39 VDD.t117 374.416
R734 VDD.t138 VDD.t49 374.416
R735 VDD.t88 VDD.t38 374.416
R736 VDD.t107 VDD.t317 374.416
R737 VDD.t278 VDD.t272 374.416
R738 VDD.t25 VDD.t318 374.416
R739 VDD.t7 VDD.t267 374.416
R740 VDD.t229 VDD.t126 374.416
R741 VDD.t79 VDD.t308 374.416
R742 VDD.t94 VDD.t334 374.416
R743 VDD.t58 VDD.t92 374.416
R744 VDD.t233 VDD.t291 318.253
R745 VDD.t199 VDD.t5 318.253
R746 VDD.t158 VDD.t218 318.253
R747 VDD.t150 VDD.t331 318.253
R748 VDD.t0 VDD.t203 318.253
R749 VDD.t262 VDD.t1 318.253
R750 VDD.t173 VDD.t211 318.253
R751 VDD.t277 VDD.t44 318.253
R752 VDD.t221 VDD.t99 318.253
R753 VDD.t293 VDD.t9 318.253
R754 VDD.t235 VDD.t298 318.253
R755 VDD.t122 VDD.t207 318.253
R756 VDD.t287 VDD.t24 318.253
R757 VDD.t304 VDD.t20 318.253
R758 VDD.t249 VDD.t127 318.253
R759 VDD.t243 VDD.t193 318.253
R760 VDD.t97 VDD.t171 318.253
R761 VDD.t333 VDD.t54 318.253
R762 VDD.t36 VDD.t101 318.253
R763 VDD.t73 VDD.t74 318.253
R764 VDD.t185 VDD.t321 318.253
R765 VDD.t270 VDD.t80 318.253
R766 VDD.t266 VDD.t43 318.253
R767 VDD.t159 VDD.t39 318.253
R768 VDD.t117 VDD.t280 318.253
R769 VDD.t256 VDD.t90 318.253
R770 VDD.t136 VDD.t138 318.253
R771 VDD.t49 VDD.t152 318.253
R772 VDD.t84 VDD.t88 318.253
R773 VDD.t38 VDD.t290 318.253
R774 VDD.t231 VDD.t247 318.253
R775 VDD.t59 VDD.t107 318.253
R776 VDD.t317 VDD.t70 318.253
R777 VDD.t167 VDD.t278 318.253
R778 VDD.t272 VDD.t312 318.253
R779 VDD.t187 VDD.t118 318.253
R780 VDD.t132 VDD.t25 318.253
R781 VDD.t318 VDD.t55 318.253
R782 VDD.t338 VDD.t7 318.253
R783 VDD.t267 VDD.t204 318.253
R784 VDD.t237 VDD.t264 318.253
R785 VDD.t177 VDD.t229 318.253
R786 VDD.t126 VDD.t213 318.253
R787 VDD.t308 VDD.t18 318.253
R788 VDD.t155 VDD.t79 318.253
R789 VDD.t225 VDD.t245 318.253
R790 VDD.t334 VDD.t14 318.253
R791 VDD.t65 VDD.t94 318.253
R792 VDD.t92 VDD.t30 318.253
R793 VDD.t29 VDD.t58 318.253
R794 VDD.n193 VDD 293.171
R795 VDD VDD.n56 288.613
R796 VDD VDD.n53 288.613
R797 VDD VDD.n49 288.613
R798 VDD VDD.n46 288.613
R799 VDD VDD.n42 288.613
R800 VDD VDD.n39 288.613
R801 VDD VDD.n35 288.613
R802 VDD VDD.n32 288.613
R803 VDD VDD.n28 288.613
R804 VDD VDD.n25 288.613
R805 VDD VDD.n21 288.613
R806 VDD VDD.n18 288.613
R807 VDD VDD.n14 288.613
R808 VDD VDD.n11 288.613
R809 VDD VDD.n7 288.613
R810 VDD VDD.n4 288.613
R811 VDD.n185 VDD 288.613
R812 VDD.n186 VDD 288.613
R813 VDD.n190 VDD 288.613
R814 VDD.t218 VDD.t68 230.889
R815 VDD.t203 VDD.t3 230.889
R816 VDD.t44 VDD.t63 230.889
R817 VDD.t9 VDD.t296 230.889
R818 VDD.t24 VDD.t273 230.889
R819 VDD.t127 VDD.t195 230.889
R820 VDD.t54 VDD.t294 230.889
R821 VDD.t74 VDD.t319 230.889
R822 VDD.t43 VDD.t169 230.889
R823 VDD.t280 VDD.t323 230.889
R824 VDD.t152 VDD.t163 230.889
R825 VDD.t290 VDD.t140 230.889
R826 VDD.t70 VDD.t47 230.889
R827 VDD.t312 VDD.t275 230.889
R828 VDD.t55 VDD.t77 230.889
R829 VDD.t204 VDD.t142 230.889
R830 VDD.t213 VDD.t285 230.889
R831 VDD.t189 VDD.t155 230.889
R832 VDD.t300 VDD.t65 230.889
R833 VDD.t209 VDD.t29 230.889
R834 VDD.t50 VDD 195.008
R835 VDD.t115 VDD 195.008
R836 VDD.t146 VDD 195.008
R837 VDD.t120 VDD 195.008
R838 VDD.t327 VDD 195.008
R839 VDD.t227 VDD 195.008
R840 VDD.t310 VDD 195.008
R841 VDD.t260 VDD 195.008
R842 VDD.t239 VDD 195.008
R843 VDD.t86 VDD 195.008
R844 VDD.t216 VDD 195.008
R845 VDD.t181 VDD 195.008
R846 VDD.t306 VDD 195.008
R847 VDD.t329 VDD 195.008
R848 VDD.t144 VDD 195.008
R849 VDD.t191 VDD 195.008
R850 VDD.t325 VDD 195.008
R851 VDD.t252 VDD 195.008
R852 VDD.t283 VDD 195.008
R853 VDD.t258 VDD 195.008
R854 VDD.t183 VDD 195.008
R855 VDD.t315 VDD 195.008
R856 VDD.t109 VDD 195.008
R857 VDD.t250 VDD 195.008
R858 VDD.t105 VDD 195.008
R859 VDD.t113 VDD 195.008
R860 VDD VDD.t241 195.008
R861 VDD VDD.t103 195.008
R862 VDD VDD.t111 195.008
R863 VDD VDD.t254 195.008
R864 VDD.t291 VDD 165.368
R865 VDD.t1 VDD 165.368
R866 VDD.t298 VDD 165.368
R867 VDD.t193 VDD 165.368
R868 VDD.t321 VDD 165.368
R869 VDD.t90 VDD 165.368
R870 VDD.t247 VDD 165.368
R871 VDD.t118 VDD 165.368
R872 VDD.t264 VDD 165.368
R873 VDD VDD.t225 165.368
R874 VDD.n204 VDD.t246 15.5636
R875 VDD.n172 VDD.t238 15.5636
R876 VDD.n158 VDD.t188 15.5636
R877 VDD.n144 VDD.t232 15.5636
R878 VDD.n130 VDD.t257 15.5636
R879 VDD.n116 VDD.t186 15.5636
R880 VDD.n102 VDD.t244 15.5636
R881 VDD.n88 VDD.t236 15.5636
R882 VDD.n74 VDD.t263 15.5636
R883 VDD.n60 VDD.t234 15.5636
R884 VDD.n195 VDD.t210 4.77854
R885 VDD.n200 VDD.t301 4.77854
R886 VDD.n181 VDD.t190 4.77854
R887 VDD.n176 VDD.t286 4.77854
R888 VDD.n167 VDD.t143 4.77854
R889 VDD.n162 VDD.t78 4.77854
R890 VDD.n153 VDD.t276 4.77854
R891 VDD.n148 VDD.t48 4.77854
R892 VDD.n139 VDD.t141 4.77854
R893 VDD.n134 VDD.t164 4.77854
R894 VDD.n125 VDD.t324 4.77854
R895 VDD.n120 VDD.t170 4.77854
R896 VDD.n111 VDD.t320 4.77854
R897 VDD.n106 VDD.t295 4.77854
R898 VDD.n97 VDD.t196 4.77854
R899 VDD.n92 VDD.t274 4.77854
R900 VDD.n83 VDD.t297 4.77854
R901 VDD.n78 VDD.t64 4.77854
R902 VDD.n69 VDD.t4 4.77854
R903 VDD.n64 VDD.t69 4.77854
R904 VDD.n198 VDD.n190 4.55932
R905 VDD.n206 VDD.n187 4.55932
R906 VDD.n186 VDD.n0 4.55932
R907 VDD.n185 VDD.n184 4.55932
R908 VDD.n170 VDD.n3 4.55932
R909 VDD.n169 VDD.n4 4.55932
R910 VDD.n164 VDD.n7 4.55932
R911 VDD.n156 VDD.n10 4.55932
R912 VDD.n155 VDD.n11 4.55932
R913 VDD.n150 VDD.n14 4.55932
R914 VDD.n142 VDD.n17 4.55932
R915 VDD.n141 VDD.n18 4.55932
R916 VDD.n136 VDD.n21 4.55932
R917 VDD.n128 VDD.n24 4.55932
R918 VDD.n127 VDD.n25 4.55932
R919 VDD.n122 VDD.n28 4.55932
R920 VDD.n114 VDD.n31 4.55932
R921 VDD.n113 VDD.n32 4.55932
R922 VDD.n108 VDD.n35 4.55932
R923 VDD.n100 VDD.n38 4.55932
R924 VDD.n99 VDD.n39 4.55932
R925 VDD.n94 VDD.n42 4.55932
R926 VDD.n86 VDD.n45 4.55932
R927 VDD.n85 VDD.n46 4.55932
R928 VDD.n80 VDD.n49 4.55932
R929 VDD.n72 VDD.n52 4.55932
R930 VDD.n71 VDD.n53 4.55932
R931 VDD.n66 VDD.n56 4.55932
R932 VDD.n197 VDD.t33 3.95308
R933 VDD.n202 VDD.t13 3.95308
R934 VDD.n183 VDD.t17 3.95308
R935 VDD.n174 VDD.t180 3.95308
R936 VDD.n165 VDD.t337 3.95308
R937 VDD.n160 VDD.t131 3.95308
R938 VDD.n151 VDD.t166 3.95308
R939 VDD.n146 VDD.t62 3.95308
R940 VDD.n137 VDD.t83 3.95308
R941 VDD.n132 VDD.t135 3.95308
R942 VDD.n123 VDD.t162 3.95308
R943 VDD.n118 VDD.t269 3.95308
R944 VDD.n109 VDD.t35 3.95308
R945 VDD.n104 VDD.t96 3.95308
R946 VDD.n95 VDD.t303 3.95308
R947 VDD.n90 VDD.t125 3.95308
R948 VDD.n81 VDD.t224 3.95308
R949 VDD.n76 VDD.t176 3.95308
R950 VDD.n67 VDD.t149 3.95308
R951 VDD.n62 VDD.t198 3.95308
R952 VDD.n203 VDD.t226 3.90058
R953 VDD.n173 VDD.t265 3.90058
R954 VDD.n159 VDD.t119 3.90058
R955 VDD.n145 VDD.t248 3.90058
R956 VDD.n131 VDD.t91 3.90058
R957 VDD.n117 VDD.t322 3.90058
R958 VDD.n103 VDD.t194 3.90058
R959 VDD.n89 VDD.t299 3.90058
R960 VDD.n75 VDD.t2 3.90058
R961 VDD.n61 VDD.t292 3.90058
R962 VDD.n205 VDD.t104 3.84351
R963 VDD.n171 VDD.t106 3.84351
R964 VDD.n157 VDD.t316 3.84351
R965 VDD.n143 VDD.t284 3.84351
R966 VDD.n129 VDD.t192 3.84351
R967 VDD.n115 VDD.t307 3.84351
R968 VDD.n101 VDD.t87 3.84351
R969 VDD.n87 VDD.t311 3.84351
R970 VDD.n73 VDD.t121 3.84351
R971 VDD.n59 VDD.t51 3.84351
R972 VDD.n192 VDD.t28 3.7805
R973 VDD.n189 VDD.t67 3.7805
R974 VDD.n179 VDD.t157 3.7805
R975 VDD.n1 VDD.t215 3.7805
R976 VDD.n5 VDD.t206 3.7805
R977 VDD.n8 VDD.t57 3.7805
R978 VDD.n12 VDD.t314 3.7805
R979 VDD.n15 VDD.t72 3.7805
R980 VDD.n19 VDD.t289 3.7805
R981 VDD.n22 VDD.t154 3.7805
R982 VDD.n26 VDD.t282 3.7805
R983 VDD.n29 VDD.t42 3.7805
R984 VDD.n33 VDD.t76 3.7805
R985 VDD.n36 VDD.t53 3.7805
R986 VDD.n40 VDD.t129 3.7805
R987 VDD.n43 VDD.t23 3.7805
R988 VDD.n47 VDD.t11 3.7805
R989 VDD.n50 VDD.t46 3.7805
R990 VDD.n54 VDD.t202 3.7805
R991 VDD.n57 VDD.t220 3.7805
R992 VDD.n194 VDD.n192 2.95854
R993 VDD.n196 VDD.n191 2.95854
R994 VDD.n199 VDD.n189 2.95854
R995 VDD.n201 VDD.n188 2.95854
R996 VDD.n180 VDD.n179 2.95854
R997 VDD.n182 VDD.n178 2.95854
R998 VDD.n177 VDD.n1 2.95854
R999 VDD.n175 VDD.n2 2.95854
R1000 VDD.n168 VDD.n5 2.95854
R1001 VDD.n166 VDD.n6 2.95854
R1002 VDD.n163 VDD.n8 2.95854
R1003 VDD.n161 VDD.n9 2.95854
R1004 VDD.n154 VDD.n12 2.95854
R1005 VDD.n152 VDD.n13 2.95854
R1006 VDD.n149 VDD.n15 2.95854
R1007 VDD.n147 VDD.n16 2.95854
R1008 VDD.n140 VDD.n19 2.95854
R1009 VDD.n138 VDD.n20 2.95854
R1010 VDD.n135 VDD.n22 2.95854
R1011 VDD.n133 VDD.n23 2.95854
R1012 VDD.n126 VDD.n26 2.95854
R1013 VDD.n124 VDD.n27 2.95854
R1014 VDD.n121 VDD.n29 2.95854
R1015 VDD.n119 VDD.n30 2.95854
R1016 VDD.n112 VDD.n33 2.95854
R1017 VDD.n110 VDD.n34 2.95854
R1018 VDD.n107 VDD.n36 2.95854
R1019 VDD.n105 VDD.n37 2.95854
R1020 VDD.n98 VDD.n40 2.95854
R1021 VDD.n96 VDD.n41 2.95854
R1022 VDD.n93 VDD.n43 2.95854
R1023 VDD.n91 VDD.n44 2.95854
R1024 VDD.n84 VDD.n47 2.95854
R1025 VDD.n82 VDD.n48 2.95854
R1026 VDD.n79 VDD.n50 2.95854
R1027 VDD.n77 VDD.n51 2.95854
R1028 VDD.n70 VDD.n54 2.95854
R1029 VDD.n68 VDD.n55 2.95854
R1030 VDD.n65 VDD.n57 2.95854
R1031 VDD.n63 VDD.n58 2.95854
R1032 VDD.n192 VDD.t255 1.53332
R1033 VDD.n189 VDD.t112 1.53332
R1034 VDD.n179 VDD.t242 1.53332
R1035 VDD.n1 VDD.t114 1.53332
R1036 VDD.n5 VDD.t251 1.53332
R1037 VDD.n8 VDD.t110 1.53332
R1038 VDD.n12 VDD.t184 1.53332
R1039 VDD.n15 VDD.t259 1.53332
R1040 VDD.n19 VDD.t253 1.53332
R1041 VDD.n22 VDD.t326 1.53332
R1042 VDD.n26 VDD.t145 1.53332
R1043 VDD.n29 VDD.t330 1.53332
R1044 VDD.n33 VDD.t182 1.53332
R1045 VDD.n36 VDD.t217 1.53332
R1046 VDD.n40 VDD.t240 1.53332
R1047 VDD.n43 VDD.t261 1.53332
R1048 VDD.n47 VDD.t228 1.53332
R1049 VDD.n50 VDD.t328 1.53332
R1050 VDD.n54 VDD.t147 1.53332
R1051 VDD.n57 VDD.t116 1.53332
R1052 VDD.n191 VDD.t31 1.31934
R1053 VDD.n191 VDD.t93 1.31934
R1054 VDD.n188 VDD.t15 1.31934
R1055 VDD.n188 VDD.t335 1.31934
R1056 VDD.n178 VDD.t19 1.31934
R1057 VDD.n178 VDD.t309 1.31934
R1058 VDD.n2 VDD.t178 1.31934
R1059 VDD.n2 VDD.t230 1.31934
R1060 VDD.n6 VDD.t339 1.31934
R1061 VDD.n6 VDD.t8 1.31934
R1062 VDD.n9 VDD.t133 1.31934
R1063 VDD.n9 VDD.t26 1.31934
R1064 VDD.n13 VDD.t168 1.31934
R1065 VDD.n13 VDD.t279 1.31934
R1066 VDD.n16 VDD.t60 1.31934
R1067 VDD.n16 VDD.t108 1.31934
R1068 VDD.n20 VDD.t85 1.31934
R1069 VDD.n20 VDD.t89 1.31934
R1070 VDD.n23 VDD.t137 1.31934
R1071 VDD.n23 VDD.t139 1.31934
R1072 VDD.n27 VDD.t160 1.31934
R1073 VDD.n27 VDD.t40 1.31934
R1074 VDD.n30 VDD.t271 1.31934
R1075 VDD.n30 VDD.t81 1.31934
R1076 VDD.n34 VDD.t37 1.31934
R1077 VDD.n34 VDD.t102 1.31934
R1078 VDD.n37 VDD.t98 1.31934
R1079 VDD.n37 VDD.t172 1.31934
R1080 VDD.n41 VDD.t305 1.31934
R1081 VDD.n41 VDD.t21 1.31934
R1082 VDD.n44 VDD.t123 1.31934
R1083 VDD.n44 VDD.t208 1.31934
R1084 VDD.n48 VDD.t222 1.31934
R1085 VDD.n48 VDD.t100 1.31934
R1086 VDD.n51 VDD.t174 1.31934
R1087 VDD.n51 VDD.t212 1.31934
R1088 VDD.n55 VDD.t151 1.31934
R1089 VDD.n55 VDD.t332 1.31934
R1090 VDD.n58 VDD.t200 1.31934
R1091 VDD.n58 VDD.t6 1.31934
R1092 VDD.n64 VDD.n63 0.3985
R1093 VDD.n69 VDD.n68 0.3985
R1094 VDD.n78 VDD.n77 0.3985
R1095 VDD.n83 VDD.n82 0.3985
R1096 VDD.n92 VDD.n91 0.3985
R1097 VDD.n97 VDD.n96 0.3985
R1098 VDD.n106 VDD.n105 0.3985
R1099 VDD.n111 VDD.n110 0.3985
R1100 VDD.n120 VDD.n119 0.3985
R1101 VDD.n125 VDD.n124 0.3985
R1102 VDD.n134 VDD.n133 0.3985
R1103 VDD.n139 VDD.n138 0.3985
R1104 VDD.n148 VDD.n147 0.3985
R1105 VDD.n153 VDD.n152 0.3985
R1106 VDD.n162 VDD.n161 0.3985
R1107 VDD.n167 VDD.n166 0.3985
R1108 VDD.n176 VDD.n175 0.3985
R1109 VDD.n182 VDD.n181 0.3985
R1110 VDD.n201 VDD.n200 0.3985
R1111 VDD.n196 VDD.n195 0.3985
R1112 VDD.n63 VDD.n62 0.3165
R1113 VDD.n68 VDD.n67 0.3165
R1114 VDD.n77 VDD.n76 0.3165
R1115 VDD.n82 VDD.n81 0.3165
R1116 VDD.n91 VDD.n90 0.3165
R1117 VDD.n96 VDD.n95 0.3165
R1118 VDD.n105 VDD.n104 0.3165
R1119 VDD.n110 VDD.n109 0.3165
R1120 VDD.n119 VDD.n118 0.3165
R1121 VDD.n124 VDD.n123 0.3165
R1122 VDD.n133 VDD.n132 0.3165
R1123 VDD.n138 VDD.n137 0.3165
R1124 VDD.n147 VDD.n146 0.3165
R1125 VDD.n152 VDD.n151 0.3165
R1126 VDD.n161 VDD.n160 0.3165
R1127 VDD.n166 VDD.n165 0.3165
R1128 VDD.n175 VDD.n174 0.3165
R1129 VDD.n183 VDD.n182 0.3165
R1130 VDD.n202 VDD.n201 0.3165
R1131 VDD.n197 VDD.n196 0.3165
R1132 VDD.n73 VDD.n72 0.2305
R1133 VDD.n87 VDD.n86 0.2305
R1134 VDD.n101 VDD.n100 0.2305
R1135 VDD.n115 VDD.n114 0.2305
R1136 VDD.n129 VDD.n128 0.2305
R1137 VDD.n143 VDD.n142 0.2305
R1138 VDD.n157 VDD.n156 0.2305
R1139 VDD.n171 VDD.n170 0.2305
R1140 VDD.n206 VDD.n205 0.2305
R1141 VDD.n65 VDD.n64 0.2125
R1142 VDD.n70 VDD.n69 0.2125
R1143 VDD.n79 VDD.n78 0.2125
R1144 VDD.n84 VDD.n83 0.2125
R1145 VDD.n93 VDD.n92 0.2125
R1146 VDD.n98 VDD.n97 0.2125
R1147 VDD.n107 VDD.n106 0.2125
R1148 VDD.n112 VDD.n111 0.2125
R1149 VDD.n121 VDD.n120 0.2125
R1150 VDD.n126 VDD.n125 0.2125
R1151 VDD.n135 VDD.n134 0.2125
R1152 VDD.n140 VDD.n139 0.2125
R1153 VDD.n149 VDD.n148 0.2125
R1154 VDD.n154 VDD.n153 0.2125
R1155 VDD.n163 VDD.n162 0.2125
R1156 VDD.n168 VDD.n167 0.2125
R1157 VDD.n177 VDD.n176 0.2125
R1158 VDD.n181 VDD.n180 0.2125
R1159 VDD.n200 VDD.n199 0.2125
R1160 VDD.n195 VDD.n194 0.2125
R1161 VDD.n66 VDD.n65 0.2085
R1162 VDD.n80 VDD.n79 0.2085
R1163 VDD.n94 VDD.n93 0.2085
R1164 VDD.n108 VDD.n107 0.2085
R1165 VDD.n122 VDD.n121 0.2085
R1166 VDD.n136 VDD.n135 0.2085
R1167 VDD.n150 VDD.n149 0.2085
R1168 VDD.n164 VDD.n163 0.2085
R1169 VDD.n184 VDD.n177 0.2085
R1170 VDD.n199 VDD.n198 0.2085
R1171 VDD.n61 VDD.n60 0.2045
R1172 VDD.n75 VDD.n74 0.2045
R1173 VDD.n89 VDD.n88 0.2045
R1174 VDD.n103 VDD.n102 0.2045
R1175 VDD.n117 VDD.n116 0.2045
R1176 VDD.n131 VDD.n130 0.2045
R1177 VDD.n145 VDD.n144 0.2045
R1178 VDD.n159 VDD.n158 0.2045
R1179 VDD.n173 VDD.n172 0.2045
R1180 VDD.n204 VDD.n203 0.2045
R1181 VDD.n71 VDD 0.1415
R1182 VDD.n85 VDD 0.1415
R1183 VDD.n99 VDD 0.1415
R1184 VDD.n113 VDD 0.1415
R1185 VDD.n127 VDD 0.1415
R1186 VDD.n141 VDD 0.1415
R1187 VDD.n155 VDD 0.1415
R1188 VDD.n169 VDD 0.1415
R1189 VDD VDD.n0 0.1415
R1190 VDD VDD.n193 0.1415
R1191 VDD.n67 VDD.n66 0.0985
R1192 VDD.n81 VDD.n80 0.0985
R1193 VDD.n95 VDD.n94 0.0985
R1194 VDD.n109 VDD.n108 0.0985
R1195 VDD.n123 VDD.n122 0.0985
R1196 VDD.n137 VDD.n136 0.0985
R1197 VDD.n151 VDD.n150 0.0985
R1198 VDD.n165 VDD.n164 0.0985
R1199 VDD.n184 VDD.n183 0.0985
R1200 VDD.n198 VDD.n197 0.0985
R1201 VDD.n60 VDD.n59 0.086
R1202 VDD.n74 VDD.n73 0.086
R1203 VDD.n88 VDD.n87 0.086
R1204 VDD.n102 VDD.n101 0.086
R1205 VDD.n116 VDD.n115 0.086
R1206 VDD.n130 VDD.n129 0.086
R1207 VDD.n144 VDD.n143 0.086
R1208 VDD.n158 VDD.n157 0.086
R1209 VDD.n172 VDD.n171 0.086
R1210 VDD.n205 VDD.n204 0.086
R1211 VDD.n62 VDD.n61 0.083
R1212 VDD.n76 VDD.n75 0.083
R1213 VDD.n90 VDD.n89 0.083
R1214 VDD.n104 VDD.n103 0.083
R1215 VDD.n118 VDD.n117 0.083
R1216 VDD.n132 VDD.n131 0.083
R1217 VDD.n146 VDD.n145 0.083
R1218 VDD.n160 VDD.n159 0.083
R1219 VDD.n174 VDD.n173 0.083
R1220 VDD.n203 VDD.n202 0.083
R1221 VDD VDD.n71 0.0775
R1222 VDD VDD.n85 0.0775
R1223 VDD VDD.n99 0.0775
R1224 VDD VDD.n113 0.0775
R1225 VDD VDD.n127 0.0775
R1226 VDD VDD.n141 0.0775
R1227 VDD VDD.n155 0.0775
R1228 VDD VDD.n169 0.0775
R1229 VDD VDD.n0 0.0775
R1230 VDD.n193 VDD 0.0775
R1231 VDD.n72 VDD 0.0755
R1232 VDD.n86 VDD 0.0755
R1233 VDD.n100 VDD 0.0755
R1234 VDD.n114 VDD 0.0755
R1235 VDD.n128 VDD 0.0755
R1236 VDD.n142 VDD 0.0755
R1237 VDD.n156 VDD 0.0755
R1238 VDD.n170 VDD 0.0755
R1239 VDD VDD.n206 0.0755
R1240 VDD VDD.n70 0.0675
R1241 VDD VDD.n84 0.0675
R1242 VDD VDD.n98 0.0675
R1243 VDD VDD.n112 0.0675
R1244 VDD VDD.n126 0.0675
R1245 VDD VDD.n140 0.0675
R1246 VDD VDD.n154 0.0675
R1247 VDD VDD.n168 0.0675
R1248 VDD.n180 VDD 0.0675
R1249 VDD.n194 VDD 0.0675
R1250 Q[4].n0 Q[4].t2 29.4195
R1251 Q[4].n2 Q[4].t3 21.1948
R1252 Q[4].n2 Q[4].t4 16.0605
R1253 Q[4].n0 Q[4].t5 11.4372
R1254 Q[4].n4 Q[4] 9.99166
R1255 Q[4] Q[4].n1 9.95
R1256 Q[4] Q[4].n5 9.14359
R1257 Q[4].n4 Q[4].n3 9.0005
R1258 Q[4].n3 Q[4].n2 8.12012
R1259 Q[4].n1 Q[4].n0 8.0005
R1260 Q[4].n5 Q[4].t0 4.5901
R1261 Q[4] Q[4].t1 3.91488
R1262 Q[4].n5 Q[4] 0.150731
R1263 Q[4] Q[4].n4 0.13775
R1264 Q[4].n1 Q[4] 0.102506
R1265 Q[4].n3 Q[4] 0.00840541
R1266 EN.n18 EN.t7 19.9538
R1267 EN.n16 EN.t11 19.9538
R1268 EN.n14 EN.t16 19.9538
R1269 EN.n12 EN.t5 19.9538
R1270 EN.n10 EN.t13 19.9538
R1271 EN.n8 EN.t0 19.9538
R1272 EN.n6 EN.t1 19.9538
R1273 EN.n4 EN.t9 19.9538
R1274 EN.n2 EN.t2 19.9538
R1275 EN.n0 EN.t8 19.9538
R1276 EN.n18 EN.t19 17.3015
R1277 EN.n16 EN.t6 17.3015
R1278 EN.n14 EN.t3 17.3015
R1279 EN.n12 EN.t15 17.3015
R1280 EN.n10 EN.t12 17.3015
R1281 EN.n8 EN.t10 17.3015
R1282 EN.n6 EN.t18 17.3015
R1283 EN.n4 EN.t14 17.3015
R1284 EN.n2 EN.t4 17.3015
R1285 EN.n0 EN.t17 17.3015
R1286 EN EN.n19 10.8498
R1287 EN.n19 EN.n18 8.0005
R1288 EN.n17 EN.n16 8.0005
R1289 EN.n15 EN.n14 8.0005
R1290 EN.n13 EN.n12 8.0005
R1291 EN.n11 EN.n10 8.0005
R1292 EN.n9 EN.n8 8.0005
R1293 EN.n7 EN.n6 8.0005
R1294 EN.n5 EN.n4 8.0005
R1295 EN.n3 EN.n2 8.0005
R1296 EN.n1 EN.n0 8.0005
R1297 EN EN.n20 6.01421
R1298 EN EN.n21 6.01421
R1299 EN EN.n22 6.01421
R1300 EN EN.n23 6.01421
R1301 EN EN.n24 6.01421
R1302 EN EN.n25 6.01421
R1303 EN EN.n26 6.01421
R1304 EN EN.n27 6.01421
R1305 EN EN.n28 6.01421
R1306 EN.n20 EN.n17 4.8361
R1307 EN.n21 EN.n15 4.8361
R1308 EN.n22 EN.n13 4.8361
R1309 EN.n23 EN.n11 4.8361
R1310 EN.n24 EN.n9 4.8361
R1311 EN.n25 EN.n7 4.8361
R1312 EN.n26 EN.n5 4.8361
R1313 EN.n27 EN.n3 4.8361
R1314 EN.n28 EN.n1 4.8361
R1315 EN.n20 EN 1.07965
R1316 EN.n21 EN 1.07965
R1317 EN.n22 EN 1.07965
R1318 EN.n23 EN 1.07965
R1319 EN.n24 EN 1.07965
R1320 EN.n25 EN 1.07965
R1321 EN.n26 EN 1.07965
R1322 EN.n27 EN 1.07965
R1323 EN.n28 EN 1.07965
R1324 EN.n19 EN 0.00742308
R1325 EN.n17 EN 0.00742308
R1326 EN.n15 EN 0.00742308
R1327 EN.n13 EN 0.00742308
R1328 EN.n11 EN 0.00742308
R1329 EN.n9 EN 0.00742308
R1330 EN.n7 EN 0.00742308
R1331 EN.n5 EN 0.00742308
R1332 EN.n3 EN 0.00742308
R1333 EN.n1 EN 0.00742308
R1334 PHI_1.n17 PHI_1.t19 26.4265
R1335 PHI_1.n15 PHI_1.t13 26.4265
R1336 PHI_1.n13 PHI_1.t2 26.4265
R1337 PHI_1.n11 PHI_1.t10 26.4265
R1338 PHI_1.n9 PHI_1.t18 26.4265
R1339 PHI_1.n7 PHI_1.t6 26.4265
R1340 PHI_1.n5 PHI_1.t9 26.4265
R1341 PHI_1.n3 PHI_1.t12 26.4265
R1342 PHI_1.n1 PHI_1.t4 26.4265
R1343 PHI_1.n0 PHI_1.t7 26.4265
R1344 PHI_1.n17 PHI_1.t16 11.7657
R1345 PHI_1.n15 PHI_1.t8 11.7657
R1346 PHI_1.n13 PHI_1.t17 11.7657
R1347 PHI_1.n11 PHI_1.t11 11.7657
R1348 PHI_1.n9 PHI_1.t5 11.7657
R1349 PHI_1.n7 PHI_1.t0 11.7657
R1350 PHI_1.n5 PHI_1.t15 11.7657
R1351 PHI_1.n3 PHI_1.t1 11.7657
R1352 PHI_1.n1 PHI_1.t3 11.7657
R1353 PHI_1.n0 PHI_1.t14 11.7657
R1354 PHI_1.n18 PHI_1 9.56151
R1355 PHI_1.n16 PHI_1 9.56151
R1356 PHI_1.n14 PHI_1 9.56151
R1357 PHI_1.n12 PHI_1 9.56151
R1358 PHI_1.n10 PHI_1 9.56151
R1359 PHI_1.n8 PHI_1 9.56151
R1360 PHI_1.n6 PHI_1 9.56151
R1361 PHI_1.n4 PHI_1 9.56151
R1362 PHI_1.n2 PHI_1 9.56151
R1363 PHI_1 PHI_1.n17 8.04713
R1364 PHI_1 PHI_1.n15 8.04713
R1365 PHI_1 PHI_1.n13 8.04713
R1366 PHI_1 PHI_1.n11 8.04713
R1367 PHI_1 PHI_1.n9 8.04713
R1368 PHI_1 PHI_1.n7 8.04713
R1369 PHI_1 PHI_1.n5 8.04713
R1370 PHI_1 PHI_1.n3 8.04713
R1371 PHI_1 PHI_1.n1 8.04713
R1372 PHI_1 PHI_1.n0 8.04713
R1373 PHI_1.n2 PHI_1 5.2583
R1374 PHI_1.n4 PHI_1 5.2583
R1375 PHI_1.n6 PHI_1 5.2583
R1376 PHI_1.n8 PHI_1 5.2583
R1377 PHI_1.n10 PHI_1 5.2583
R1378 PHI_1.n12 PHI_1 5.2583
R1379 PHI_1.n14 PHI_1 5.2583
R1380 PHI_1.n16 PHI_1 5.2583
R1381 PHI_1 PHI_1.n18 5.2583
R1382 PHI_1 PHI_1.n2 0.3587
R1383 PHI_1 PHI_1.n4 0.3587
R1384 PHI_1 PHI_1.n6 0.3587
R1385 PHI_1 PHI_1.n8 0.3587
R1386 PHI_1 PHI_1.n10 0.3587
R1387 PHI_1 PHI_1.n12 0.3587
R1388 PHI_1 PHI_1.n14 0.3587
R1389 PHI_1 PHI_1.n16 0.3587
R1390 PHI_1.n18 PHI_1 0.3587
R1391 PHI_2.n17 PHI_2.t6 26.4265
R1392 PHI_2.n15 PHI_2.t7 26.4265
R1393 PHI_2.n13 PHI_2.t5 26.4265
R1394 PHI_2.n11 PHI_2.t12 26.4265
R1395 PHI_2.n9 PHI_2.t14 26.4265
R1396 PHI_2.n7 PHI_2.t16 26.4265
R1397 PHI_2.n5 PHI_2.t10 26.4265
R1398 PHI_2.n3 PHI_2.t13 26.4265
R1399 PHI_2.n1 PHI_2.t15 26.4265
R1400 PHI_2.n0 PHI_2.t4 26.4265
R1401 PHI_2.n17 PHI_2.t0 11.7657
R1402 PHI_2.n15 PHI_2.t8 11.7657
R1403 PHI_2.n13 PHI_2.t2 11.7657
R1404 PHI_2.n11 PHI_2.t17 11.7657
R1405 PHI_2.n9 PHI_2.t11 11.7657
R1406 PHI_2.n7 PHI_2.t19 11.7657
R1407 PHI_2.n5 PHI_2.t1 11.7657
R1408 PHI_2.n3 PHI_2.t9 11.7657
R1409 PHI_2.n1 PHI_2.t3 11.7657
R1410 PHI_2.n0 PHI_2.t18 11.7657
R1411 PHI_2.n18 PHI_2 9.23499
R1412 PHI_2.n16 PHI_2 9.23499
R1413 PHI_2.n14 PHI_2 9.23499
R1414 PHI_2.n12 PHI_2 9.23499
R1415 PHI_2.n10 PHI_2 9.23499
R1416 PHI_2.n8 PHI_2 9.23499
R1417 PHI_2.n6 PHI_2 9.23499
R1418 PHI_2.n4 PHI_2 9.23499
R1419 PHI_2.n2 PHI_2 9.23499
R1420 PHI_2 PHI_2.n17 8.04257
R1421 PHI_2 PHI_2.n15 8.04257
R1422 PHI_2 PHI_2.n13 8.04257
R1423 PHI_2 PHI_2.n11 8.04257
R1424 PHI_2 PHI_2.n9 8.04257
R1425 PHI_2 PHI_2.n7 8.04257
R1426 PHI_2 PHI_2.n5 8.04257
R1427 PHI_2 PHI_2.n3 8.04257
R1428 PHI_2 PHI_2.n1 8.04257
R1429 PHI_2 PHI_2.n0 8.04257
R1430 PHI_2.n2 PHI_2 3.0407
R1431 PHI_2.n4 PHI_2 3.0407
R1432 PHI_2.n6 PHI_2 3.0407
R1433 PHI_2.n8 PHI_2 3.0407
R1434 PHI_2.n10 PHI_2 3.0407
R1435 PHI_2.n12 PHI_2 3.0407
R1436 PHI_2.n14 PHI_2 3.0407
R1437 PHI_2.n16 PHI_2 3.0407
R1438 PHI_2.n18 PHI_2 3.0407
R1439 PHI_2 PHI_2.n2 2.5763
R1440 PHI_2 PHI_2.n4 2.5763
R1441 PHI_2 PHI_2.n6 2.5763
R1442 PHI_2 PHI_2.n8 2.5763
R1443 PHI_2 PHI_2.n10 2.5763
R1444 PHI_2 PHI_2.n12 2.5763
R1445 PHI_2 PHI_2.n14 2.5763
R1446 PHI_2 PHI_2.n16 2.5763
R1447 PHI_2 PHI_2.n18 2.5763
R1448 Q[6].n0 Q[6].t2 29.4195
R1449 Q[6].n2 Q[6].t5 21.1948
R1450 Q[6].n2 Q[6].t3 16.0605
R1451 Q[6].n0 Q[6].t4 11.4372
R1452 Q[6].n4 Q[6] 9.99166
R1453 Q[6] Q[6].n1 9.95
R1454 Q[6] Q[6].n5 9.14359
R1455 Q[6].n4 Q[6].n3 9.0005
R1456 Q[6].n3 Q[6].n2 8.12012
R1457 Q[6].n1 Q[6].n0 8.0005
R1458 Q[6].n5 Q[6].t0 4.5901
R1459 Q[6] Q[6].t1 3.91488
R1460 Q[6].n5 Q[6] 0.150731
R1461 Q[6] Q[6].n4 0.13775
R1462 Q[6].n1 Q[6] 0.102506
R1463 Q[6].n3 Q[6] 0.00840541
R1464 gc[2] gc[2].n0 16.6226
R1465 gc[2].n0 gc[2].t0 4.57685
R1466 gc[2] gc[2].t1 4.33791
R1467 gc[2].n0 gc[2] 0.0122931
R1468 gc[8] gc[8].n0 16.6476
R1469 gc[8].n0 gc[8].t0 4.57685
R1470 gc[8] gc[8].t1 4.33791
R1471 gc[8].n0 gc[8] 0.0122931
R1472 D_in.n0 D_in.t1 29.4195
R1473 D_in.n0 D_in.t0 11.4372
R1474 D_in D_in.n1 9.95
R1475 D_in.n1 D_in.n0 8.0005
R1476 D_in.n1 D_in 0.102506
R1477 Q[2].n0 Q[2].t2 29.4195
R1478 Q[2].n2 Q[2].t4 21.1948
R1479 Q[2].n2 Q[2].t5 16.0605
R1480 Q[2].n0 Q[2].t3 11.4372
R1481 Q[2].n4 Q[2] 9.99166
R1482 Q[2] Q[2].n1 9.95
R1483 Q[2] Q[2].n5 9.16834
R1484 Q[2].n4 Q[2].n3 9.0005
R1485 Q[2].n3 Q[2].n2 8.12012
R1486 Q[2].n1 Q[2].n0 8.0005
R1487 Q[2].n5 Q[2].t0 4.5901
R1488 Q[2] Q[2].t1 3.91488
R1489 Q[2].n5 Q[2] 0.150731
R1490 Q[2] Q[2].n4 0.13775
R1491 Q[2].n1 Q[2] 0.102506
R1492 Q[2].n3 Q[2] 0.00840541
R1493 Q[7].n0 Q[7].t4 29.4195
R1494 Q[7].n2 Q[7].t5 21.1948
R1495 Q[7].n2 Q[7].t3 16.0605
R1496 Q[7].n0 Q[7].t2 11.4372
R1497 Q[7].n4 Q[7] 9.99166
R1498 Q[7] Q[7].n1 9.95
R1499 Q[7] Q[7].n5 9.14359
R1500 Q[7].n4 Q[7].n3 9.0005
R1501 Q[7].n3 Q[7].n2 8.12012
R1502 Q[7].n1 Q[7].n0 8.0005
R1503 Q[7].n5 Q[7].t0 4.5901
R1504 Q[7] Q[7].t1 3.91488
R1505 Q[7].n5 Q[7] 0.150731
R1506 Q[7] Q[7].n4 0.13775
R1507 Q[7].n1 Q[7] 0.102506
R1508 Q[7].n3 Q[7] 0.00840541
R1509 gc[5] gc[5].n0 16.6626
R1510 gc[5].n0 gc[5].t0 4.57685
R1511 gc[5] gc[5].t1 4.33791
R1512 gc[5].n0 gc[5] 0.0122931
R1513 Q[1].n0 Q[1].t4 29.4195
R1514 Q[1].n2 Q[1].t5 21.1948
R1515 Q[1].n2 Q[1].t3 16.0605
R1516 Q[1].n0 Q[1].t2 11.4372
R1517 Q[1].n4 Q[1] 9.99166
R1518 Q[1] Q[1].n1 9.95
R1519 Q[1] Q[1].n5 9.06259
R1520 Q[1].n4 Q[1].n3 9.0005
R1521 Q[1].n3 Q[1].n2 8.12012
R1522 Q[1].n1 Q[1].n0 8.0005
R1523 Q[1].n5 Q[1].t0 4.5901
R1524 Q[1] Q[1].t1 3.91488
R1525 Q[1].n5 Q[1] 0.150731
R1526 Q[1] Q[1].n4 0.13775
R1527 Q[1].n1 Q[1] 0.102506
R1528 Q[1].n3 Q[1] 0.00840541
R1529 gc[7] gc[7].n0 16.6126
R1530 gc[7].n0 gc[7].t0 4.57685
R1531 gc[7] gc[7].t1 4.33791
R1532 gc[7].n0 gc[7] 0.0122931
R1533 Q[10].n0 Q[10].t2 21.1948
R1534 Q[10].n0 Q[10].t3 16.0605
R1535 Q[10] Q[10].n2 9.16609
R1536 Q[10] Q[10].n1 9.13775
R1537 Q[10].n1 Q[10].n0 8.12012
R1538 Q[10].n2 Q[10].t0 4.5901
R1539 Q[10] Q[10].t1 3.91488
R1540 Q[10].n2 Q[10] 0.150731
R1541 Q[10].n1 Q[10] 0.00840541
R1542 gc[1] gc[1].n0 16.6451
R1543 gc[1].n0 gc[1].t0 4.57685
R1544 gc[1] gc[1].t1 4.33791
R1545 gc[1].n0 gc[1] 0.0122931
R1546 Q[3].n0 Q[3].t5 29.4195
R1547 Q[3].n2 Q[3].t4 21.1948
R1548 Q[3].n2 Q[3].t3 16.0605
R1549 Q[3].n0 Q[3].t2 11.4372
R1550 Q[3].n4 Q[3] 9.99166
R1551 Q[3] Q[3].n1 9.95
R1552 Q[3] Q[3].n5 9.14584
R1553 Q[3].n4 Q[3].n3 9.0005
R1554 Q[3].n3 Q[3].n2 8.12012
R1555 Q[3].n1 Q[3].n0 8.0005
R1556 Q[3].n5 Q[3].t0 4.5901
R1557 Q[3] Q[3].t1 3.91488
R1558 Q[3].n5 Q[3] 0.150731
R1559 Q[3] Q[3].n4 0.13775
R1560 Q[3].n1 Q[3] 0.102506
R1561 Q[3].n3 Q[3] 0.00840541
R1562 Q[5].n0 Q[5].t2 29.4195
R1563 Q[5].n2 Q[5].t3 21.1948
R1564 Q[5].n2 Q[5].t5 16.0605
R1565 Q[5].n0 Q[5].t4 11.4372
R1566 Q[5].n4 Q[5] 9.99166
R1567 Q[5] Q[5].n1 9.95
R1568 Q[5] Q[5].n5 9.14359
R1569 Q[5].n4 Q[5].n3 9.0005
R1570 Q[5].n3 Q[5].n2 8.12012
R1571 Q[5].n1 Q[5].n0 8.0005
R1572 Q[5].n5 Q[5].t0 4.5901
R1573 Q[5] Q[5].t1 3.91488
R1574 Q[5].n5 Q[5] 0.150731
R1575 Q[5] Q[5].n4 0.13775
R1576 Q[5].n1 Q[5] 0.102506
R1577 Q[5].n3 Q[5] 0.00840541
R1578 Q[9].n0 Q[9].t4 29.4195
R1579 Q[9].n2 Q[9].t3 21.1948
R1580 Q[9].n2 Q[9].t5 16.0605
R1581 Q[9].n0 Q[9].t2 11.4372
R1582 Q[9].n4 Q[9] 9.99166
R1583 Q[9] Q[9].n1 9.95
R1584 Q[9] Q[9].n5 9.14359
R1585 Q[9].n4 Q[9].n3 9.0005
R1586 Q[9].n3 Q[9].n2 8.12012
R1587 Q[9].n1 Q[9].n0 8.0005
R1588 Q[9].n5 Q[9].t0 4.5901
R1589 Q[9] Q[9].t1 3.91488
R1590 Q[9].n5 Q[9] 0.150731
R1591 Q[9] Q[9].n4 0.13775
R1592 Q[9].n1 Q[9] 0.102506
R1593 Q[9].n3 Q[9] 0.00840541
R1594 Q[8].n0 Q[8].t3 29.4195
R1595 Q[8].n2 Q[8].t4 21.1948
R1596 Q[8].n2 Q[8].t5 16.0605
R1597 Q[8].n0 Q[8].t2 11.4372
R1598 Q[8].n4 Q[8] 9.99166
R1599 Q[8] Q[8].n1 9.95
R1600 Q[8] Q[8].n5 9.14359
R1601 Q[8].n4 Q[8].n3 9.0005
R1602 Q[8].n3 Q[8].n2 8.12012
R1603 Q[8].n1 Q[8].n0 8.0005
R1604 Q[8].n5 Q[8].t0 4.5901
R1605 Q[8] Q[8].t1 3.91488
R1606 Q[8].n5 Q[8] 0.150731
R1607 Q[8] Q[8].n4 0.13775
R1608 Q[8].n1 Q[8] 0.102506
R1609 Q[8].n3 Q[8] 0.00840541
R1610 gc[4] gc[4].n0 16.6314
R1611 gc[4].n0 gc[4].t0 4.57685
R1612 gc[4] gc[4].t1 4.33791
R1613 gc[4].n0 gc[4] 0.0122931
R1614 gc[9] gc[9].n0 16.6301
R1615 gc[9].n0 gc[9].t0 4.57685
R1616 gc[9] gc[9].t1 4.33791
R1617 gc[9].n0 gc[9] 0.0122931
R1618 gc[3] gc[3].n0 16.6089
R1619 gc[3].n0 gc[3].t0 4.57685
R1620 gc[3] gc[3].t1 4.33791
R1621 gc[3].n0 gc[3] 0.0122931
R1622 gc[6] gc[6].n0 16.6401
R1623 gc[6].n0 gc[6].t0 4.57685
R1624 gc[6] gc[6].t1 4.33791
R1625 gc[6].n0 gc[6] 0.0122931
R1626 gc[10] gc[10].n0 16.6539
R1627 gc[10].n0 gc[10].t0 4.57685
R1628 gc[10] gc[10].t1 4.33791
R1629 gc[10].n0 gc[10] 0.0122931
C0 EN a_48974_158# 0.11055f
C1 PHI_2 a_48826_158# 0
C2 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_39302_38# 0.00242f
C3 PHI_2 a_42586_n387# 0
C4 gc[8] a_42978_n387# 0
C5 a_17626_158# EN 0.00101f
C6 a_n1462_n384# PHI_2 0.03321f
C7 Q[5] a_26478_158# 0.11433f
C8 a_24358_38# a_24014_158# 0.57845f
C9 a_23498_n384# a_25494_n402# 0
C10 a_58022_38# gc[10] 0.01014f
C11 a_5294_158# a_6774_n402# 0.00268f
C12 PHI_1 a_50454_n402# 0.01733f
C13 EN Q[9] 0.513f
C14 a_17774_158# PHI_2 0.04895f
C15 a_38442_n384# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C16 a_17978_158# PHI_1 0.00534f
C17 EN a_45542_38# 0.0522f
C18 gc[7] a_38810_n387# 0
C19 a_11878_38# Q[2] 0.00242f
C20 gc[7] a_38442_n384# 0.00668f
C21 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_1862_38# 0.00242f
C22 a_18018_n387# a_18118_38# 0
C23 a_n1094_158# PHI_1 0.00201f
C24 PHI_2 a_46663_n425# 0
C25 a_5146_158# PHI_2 0
C26 gc[8] a_45050_n387# 0
C27 EN a_42734_158# 0.11055f
C28 a_8102_38# VDD 0.32599f
C29 a_2983_n425# Q[1] 0.00241f
C30 a_17258_n384# PHI_2 0.03321f
C31 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[9] 0.23535f
C32 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_11878_38# 0.2556f
C33 a_20238_158# EN 0.11443f
C34 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_n1930_n402# 0.00116f
C35 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_38810_n387# 0
C36 PHI_1 a_44214_n402# 0.01733f
C37 EN a_47990_n402# 0.08752f
C38 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_38442_n384# 0.36162f
C39 gc[8] a_45402_158# 0
C40 a_5498_158# EN 0.00368f
C41 PHI_2 a_42978_n387# 0
C42 a_18018_n387# a_17774_158# 0.01595f
C43 PHI_1 a_48974_158# 0.01882f
C44 a_57162_n384# gc[10] 0.00668f
C45 a_24358_38# a_23030_n402# 0.02403f
C46 a_23498_n384# a_24014_158# 0.30053f
C47 a_14342_38# gc[3] 0.01014f
C48 a_17626_158# PHI_1 0.00201f
C49 a_38958_158# DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C50 a_16790_n402# PHI_2 0.02762f
C51 a_11018_n384# Q[2] 0.36203f
C52 gc[7] a_39202_n387# 0
C53 EN a_44682_n384# 0.05124f
C54 Q[9] PHI_1 0.05798f
C55 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_1002_n384# 0.36162f
C56 a_50454_n402# a_51782_38# 0.02403f
C57 gc[7] a_38958_158# 0.01553f
C58 gc[2] a_7962_158# 0
C59 PHI_1 a_45542_38# 0.01261f
C60 gc[3] Q[2] 0.17162f
C61 a_n946_158# a_534_n402# 0.00268f
C62 EN a_41750_n402# 0.08752f
C63 gc[8] a_45442_n387# 0
C64 PHI_2 a_45050_n387# 0
C65 a_7242_n384# VDD 0.42245f
C66 a_19254_n402# PHI_2 0.60119f
C67 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_11018_n384# 0
C68 a_11738_158# VDD 0.01506f
C69 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_50922_n384# 0
C70 PHI_2 a_7962_158# 0.00422f
C71 PHI_1 a_42734_158# 0.01882f
C72 a_2983_n425# PHI_2 0
C73 PHI_2 a_45402_158# 0.00422f
C74 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_38958_158# 0.01536f
C75 a_13014_n402# a_14342_38# 0.02403f
C76 a_7610_n387# a_7242_n384# 0.00194f
C77 a_8002_n387# a_8102_38# 0
C78 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_19722_n384# 0
C79 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[3] 0.23535f
C80 Q[8] VDD 0.56326f
C81 a_20238_158# PHI_1 0.01804f
C82 a_58022_38# Q[10] 0.25874f
C83 Q[7] a_39302_38# 0.25874f
C84 PHI_1 a_47990_n402# 0.70141f
C85 a_23498_n384# a_23030_n402# 0.30528f
C86 a_57678_158# gc[10] 0.01553f
C87 a_5498_158# PHI_1 0.00534f
C88 a_13482_n384# gc[3] 0.00668f
C89 EN a_45198_158# 0.11443f
C90 EN a_36738_n387# 0.00577f
C91 a_50454_n402# a_50922_n384# 0.30528f
C92 a_1518_158# EN 0.11443f
C93 a_11878_38# VDD 0.32599f
C94 PHI_1 a_44682_n384# 0.01277f
C95 PHI_2 a_58022_38# 0.03174f
C96 Q[9] a_51782_38# 0.25874f
C97 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD 0.34237f
C98 PHI_2 a_45442_n387# 0
C99 a_24358_38# EN 0.05124f
C100 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_13014_n402# 0.16689f
C101 a_26822_38# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00242f
C102 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_51438_158# 0.00144f
C103 PHI_1 a_41750_n402# 0.70141f
C104 a_7242_n384# a_8102_38# 0.00888f
C105 a_7758_158# a_7610_158# 0
C106 a_13014_n402# a_13482_n384# 0.30528f
C107 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_13850_n387# 0
C108 PHI_2 a_45050_158# 0
C109 a_1370_n387# PHI_2 0
C110 a_57162_n384# Q[10] 0.00101f
C111 a_5146_158# a_5294_158# 0
C112 Q[7] a_38442_n384# 0.00101f
C113 a_14242_n387# a_14342_38# 0
C114 a_13850_n387# a_13482_n384# 0.00194f
C115 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gc[4] 0.33472f
C116 a_1862_38# Q[1] 0.25874f
C117 a_11534_158# Q[2] 0.01552f
C118 a_20582_38# a_20238_158# 0.57845f
C119 gc[7] a_36346_n387# 0
C120 EN a_39162_158# 0.00368f
C121 a_50454_n402# a_51438_158# 0.07055f
C122 VDD DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42635f
C123 VDD a_26822_38# 0.32599f
C124 a_11018_n384# VDD 0.4225f
C125 PHI_1 a_45198_158# 0.01804f
C126 PHI_2 a_57162_n384# 0.07395f
C127 PHI_2 a_49178_158# 0.00411f
C128 a_1518_158# PHI_1 0.01804f
C129 gc[7] VDD 0.26766f
C130 Q[9] a_50922_n384# 0.00101f
C131 gc[3] VDD 0.26766f
C132 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[1] 0.23535f
C133 a_23498_n384# EN 0.05108f
C134 gc[5] a_23866_n387# 0
C135 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_11534_158# 0.09501f
C136 a_20482_n387# PHI_2 0
C137 a_17978_158# gc[4] 0
C138 VDD DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42635f
C139 a_n946_158# a_n1094_158# 0
C140 a_534_n402# a_n602_38# 0
C141 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_40423_n425# 0.0097f
C142 a_14342_38# Q[3] 0.25874f
C143 a_1762_n387# PHI_2 0
C144 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_20090_n387# 0
C145 a_24358_38# PHI_1 0.01314f
C146 gc[7] a_40423_n425# 0.00113f
C147 PHI_2 a_39302_38# 0.03174f
C148 a_57678_158# Q[10] 0.11433f
C149 Q[7] a_38958_158# 0.11433f
C150 gc[6] EN 0.44384f
C151 VDD DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C152 VDD DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C153 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD 0.34237f
C154 a_1002_n384# Q[1] 0.00101f
C155 a_49318_38# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.2556f
C156 EN a_38810_158# 0.00101f
C157 a_5498_158# a_5638_38# 0.00109f
C158 a_19722_n384# a_20238_158# 0.30053f
C159 a_1862_38# PHI_2 0.03174f
C160 a_13014_n402# VDD 1.03607f
C161 PHI_1 a_39162_158# 0.00477f
C162 PHI_2 a_57678_158# 0.04011f
C163 Q[9] a_51438_158# 0.11433f
C164 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[3] 0.01102f
C165 gc[5] a_24258_n387# 0
C166 a_11738_158# a_11878_38# 0.00109f
C167 a_24218_158# PHI_2 0.00411f
C168 a_49178_158# gc[9] 0
C169 VDD a_29738_n384# 0.4225f
C170 a_13482_n384# Q[3] 0.00101f
C171 a_534_n402# a_n1462_n384# 0
C172 PHI_2 a_n1930_n402# 0.02723f
C173 a_25494_n402# gc[5] 0.00985f
C174 EN a_43078_38# 0.05124f
C175 PHI_2 a_38810_n387# 0
C176 a_23498_n384# PHI_1 0.0533f
C177 a_14202_158# EN 0.00368f
C178 PHI_2 a_38442_n384# 0.07395f
C179 a_30598_38# gc[6] 0.00972f
C180 a_48458_n384# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C181 a_1370_158# PHI_2 0
C182 EN DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C183 gc[6] PHI_1 0.01023f
C184 a_1002_n384# PHI_2 0.07395f
C185 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[1] 0.08575f
C186 a_11534_158# VDD 0.56047f
C187 a_20238_158# gc[4] 0.01553f
C188 a_39302_38# a_37974_n402# 0.02403f
C189 PHI_1 a_38810_158# 0.00164f
C190 a_48458_n384# a_48826_158# 0.00294f
C191 a_1722_158# EN 0.00368f
C192 Q[4] DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C193 VDD gc[10] 0.26726f
C194 a_14342_38# PHI_2 0.03174f
C195 a_23866_158# PHI_2 0
C196 gc[5] a_26682_158# 0
C197 VDD a_31734_n402# 1.03607f
C198 a_26330_n387# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C199 gc[2] Q[2] 0.22418f
C200 a_24014_158# gc[5] 0.01329f
C201 gc[8] a_42938_158# 0
C202 PHI_2 a_39202_n387# 0
C203 EN a_42218_n384# 0.05108f
C204 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_56694_n402# 0
C205 a_13850_158# EN 0.00101f
C206 a_11738_158# gc[3] 0
C207 PHI_2 a_38958_158# 0.04011f
C208 Q[2] PHI_2 0.63578f
C209 PHI_1 a_43078_38# 0.01314f
C210 a_14202_158# PHI_1 0.00477f
C211 Q[7] VDD 0.56326f
C212 a_50454_n402# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.16689f
C213 Q[4] VDD 0.56326f
C214 EN a_5146_n387# 0.0022f
C215 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_44214_n402# 0
C216 Q[3] VDD 0.56326f
C217 VDD a_55558_38# 0.32599f
C218 a_11018_n384# a_11878_38# 0.00888f
C219 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_2 0.45413f
C220 a_18118_38# a_17978_158# 0.00109f
C221 gc[1] Q[1] 0.22418f
C222 a_38442_n384# a_37974_n402# 0.30528f
C223 PHI_1 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C224 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C225 Q[4] a_21703_n425# 0.00241f
C226 Q[7] a_40423_n425# 0.00241f
C227 Q[8] DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01102f
C228 a_13482_n384# PHI_2 0.07395f
C229 a_59143_n425# gc[10] 0.00113f
C230 a_11878_38# gc[3] 0.00972f
C231 Q[6] EN 0.513f
C232 VDD a_30254_158# 0.56047f
C233 a_23030_n402# gc[5] 0.00985f
C234 a_1722_158# PHI_1 0.00477f
C235 PHI_2 a_42938_158# 0.00411f
C236 a_24014_158# a_23866_n387# 0
C237 a_17978_158# a_17774_158# 0.01151f
C238 Q[1] VDD 0.56326f
C239 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[2] 0.01102f
C240 a_n1462_n384# a_n1094_158# 0.00294f
C241 PHI_1 a_42218_n384# 0.0533f
C242 a_13850_158# PHI_1 0.00164f
C243 gc[8] VDD 0.26766f
C244 gc[6] Q[5] 0.17162f
C245 a_48974_158# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.09501f
C246 a_9223_n425# gc[2] 0.00113f
C247 EN a_5538_n387# 0.00577f
C248 VDD a_54698_n384# 0.4225f
C249 a_7758_158# EN 0.11443f
C250 a_9223_n425# PHI_2 0
C251 a_13014_n402# a_11878_38# 0
C252 gc[2] gc[1] 0.01049f
C253 PHI_2 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C254 a_38958_158# a_37974_n402# 0.07055f
C255 Q[9] DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01102f
C256 a_48974_158# a_48826_158# 0
C257 gc[7] DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.33472f
C258 a_47990_n402# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C259 a_55214_158# a_56694_n402# 0.00268f
C260 a_n1094_n387# PHI_2 0
C261 a_57530_n387# gc[10] 0
C262 gc[1] PHI_2 0.31085f
C263 VDD Q[10] 0.38176f
C264 a_11018_n384# gc[3] 0.00668f
C265 a_11738_158# a_11534_158# 0.01151f
C266 VDD a_36838_38# 0.32599f
C267 VDD a_29270_n402# 1.00028f
C268 PHI_2 a_42586_158# 0
C269 a_15463_n425# gc[3] 0.00113f
C270 PHI_2 a_36346_n387# 0
C271 a_24014_158# a_24258_n387# 0.01595f
C272 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_19254_n402# 0
C273 a_17626_158# a_17774_158# 0
C274 a_55066_n387# a_55214_158# 0
C275 Q[6] PHI_1 0.05798f
C276 gc[2] VDD 0.26766f
C277 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_44682_n384# 0
C278 a_24014_158# a_25494_n402# 0.00268f
C279 VDD a_36698_158# 0.01506f
C280 PHI_2 VDD 4.64303f
C281 a_47990_n402# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00116f
C282 a_49318_38# a_49178_158# 0.00109f
C283 a_7610_n387# gc[2] 0
C284 a_42586_n387# a_42734_158# 0
C285 gc[7] DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.23535f
C286 a_36346_n387# a_35978_n384# 0.00194f
C287 a_23498_n384# gc[4] 0
C288 a_11534_158# a_11878_38# 0.57845f
C289 a_30458_158# VDD 0.01506f
C290 gc[5] EN 0.44384f
C291 a_13014_n402# a_11018_n384# 0
C292 a_7610_n387# PHI_2 0
C293 a_17258_n384# a_17626_158# 0.00294f
C294 PHI_2 a_21703_n425# 0
C295 a_7758_158# PHI_1 0.01804f
C296 a_54230_n402# a_56694_n402# 0
C297 PHI_2 a_40423_n425# 0
C298 a_n702_n387# PHI_2 0
C299 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_56694_n402# 0.16689f
C300 a_57922_n387# gc[10] 0
C301 VDD DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42635f
C302 a_13014_n402# gc[3] 0.00985f
C303 a_59143_n425# Q[10] 0.00241f
C304 VDD a_35978_n384# 0.4225f
C305 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD 0.34237f
C306 a_13850_n387# gc[3] 0
C307 a_55458_n387# a_55214_158# 0.01595f
C308 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_45198_158# 0.00144f
C309 a_23030_n402# a_25494_n402# 0
C310 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN 0.65271f
C311 PHI_2 a_59143_n425# 0
C312 a_1862_38# a_534_n402# 0.02403f
C313 a_8102_38# gc[2] 0.01014f
C314 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD 0.34237f
C315 a_8002_n387# gc[2] 0
C316 a_42978_n387# a_42734_158# 0.01595f
C317 VDD gc[9] 0.26766f
C318 a_8102_38# PHI_2 0.03174f
C319 a_11534_158# a_11018_n384# 0.30053f
C320 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[4] 0.01102f
C321 a_7610_n387# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C322 a_8002_n387# PHI_2 0
C323 a_30106_158# VDD 0.00491f
C324 PHI_2 a_20090_n387# 0
C325 EN a_23866_n387# 0.0022f
C326 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[3] 0.01068f
C327 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_55214_158# 0.09501f
C328 a_54230_n402# a_55214_158# 0.07055f
C329 a_534_n402# a_n1930_n402# 0
C330 gc[5] PHI_1 0.01023f
C331 a_11534_158# gc[3] 0.01329f
C332 a_7610_158# EN 0.00101f
C333 gc[8] Q[8] 0.22418f
C334 VDD a_37974_n402# 1.03607f
C335 EN DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C336 a_14242_n387# gc[3] 0
C337 a_23030_n402# a_24014_158# 0.07055f
C338 a_n742_158# EN 0.00368f
C339 a_45402_158# a_45542_38# 0.00109f
C340 VDD a_51642_158# 0.01506f
C341 a_20442_158# VDD 0.01506f
C342 a_11386_n387# EN 0.0022f
C343 Q[7] DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C344 a_1002_n384# a_534_n402# 0.30528f
C345 PHI_2 a_57530_n387# 0
C346 a_7242_n384# gc[2] 0.00668f
C347 a_20238_158# a_19254_n402# 0.07055f
C348 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C349 a_7242_n384# PHI_2 0.07395f
C350 a_36346_n387# a_36494_158# 0
C351 a_11534_158# a_13014_n402# 0.00268f
C352 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_8102_38# 0.00242f
C353 a_11738_158# PHI_2 0.00411f
C354 EN a_56694_n402# 0.08694f
C355 Q[7] gc[7] 0.22418f
C356 a_15463_n425# Q[3] 0.00241f
C357 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_10550_n402# 0
C358 EN a_24258_n387# 0.00577f
C359 Q[3] gc[3] 0.22418f
C360 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_54230_n402# 0.00116f
C361 VDD a_5294_158# 0.56047f
C362 a_25494_n402# EN 0.08694f
C363 a_45050_n387# a_44682_n384# 0.00194f
C364 a_45442_n387# a_45542_38# 0
C365 Q[8] PHI_2 0.63578f
C366 a_5538_n387# a_5638_38# 0
C367 VDD a_36494_158# 0.56047f
C368 a_5146_n387# a_4778_n384# 0.00194f
C369 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_6774_n402# 0
C370 a_33062_38# VDD 0.32599f
C371 EN a_55066_n387# 0.0022f
C372 Q[7] DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01102f
C373 a_7610_158# PHI_1 0.00164f
C374 Q[7] DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C375 a_20090_158# VDD 0.00491f
C376 VDD a_51290_158# 0.00491f
C377 PHI_1 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.01636f
C378 a_11778_n387# EN 0.00577f
C379 a_31734_n402# a_29738_n384# 0
C380 EN a_4310_n402# 0.08752f
C381 a_11878_38# PHI_2 0.03207f
C382 PHI_2 a_57922_n387# 0
C383 a_n742_158# PHI_1 0.00534f
C384 a_48974_158# a_49178_158# 0.01151f
C385 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_25962_n384# 0.36162f
C386 a_13014_n402# Q[3] 0.00225f
C387 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_2 0.45413f
C388 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_534_n402# 0
C389 gc[8] gc[7] 0.01049f
C390 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_7242_n384# 0.36162f
C391 a_26722_n387# a_26822_38# 0
C392 EN a_55214_158# 0.11055f
C393 EN a_26682_158# 0.00368f
C394 a_11386_158# EN 0.00101f
C395 gc[5] Q[5] 0.22418f
C396 a_24014_158# EN 0.11055f
C397 VDD a_32922_158# 0.01506f
C398 a_55214_158# a_55418_158# 0.01151f
C399 PHI_1 a_56694_n402# 0.01733f
C400 a_45050_n387# a_45198_158# 0
C401 VDD a_35510_n402# 1.00028f
C402 EN a_55458_n387# 0.00577f
C403 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[1] 0.01102f
C404 a_32202_n384# VDD 0.42245f
C405 a_13998_158# a_14342_38# 0.57845f
C406 Q[8] gc[9] 0.17162f
C407 gc[8] DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.23535f
C408 a_25494_n402# PHI_1 0.01733f
C409 gc[7] a_36838_38# 0.00972f
C410 VDD a_25962_n384# 0.42245f
C411 a_11018_n384# gc[2] 0
C412 a_45402_158# a_45198_158# 0.01151f
C413 a_45050_158# a_44682_n384# 0.00294f
C414 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_29270_n402# 0
C415 a_30254_158# a_29738_n384# 0.30053f
C416 PHI_2 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C417 PHI_2 a_26822_38# 0.03174f
C418 a_11018_n384# PHI_2 0.03321f
C419 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_26478_158# 0.01536f
C420 gc[7] a_36698_158# 0
C421 gc[2] gc[3] 0.01049f
C422 a_20482_n387# a_20238_158# 0.01595f
C423 gc[7] PHI_2 0.31085f
C424 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_36838_38# 0.2556f
C425 a_15463_n425# PHI_2 0
C426 PHI_1 a_4310_n402# 0.70141f
C427 gc[3] PHI_2 0.31085f
C428 EN DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C429 EN a_54230_n402# 0.08752f
C430 EN a_51290_n387# 0.0022f
C431 Q[8] a_48826_n387# 0
C432 EN a_26330_158# 0.00101f
C433 a_534_n402# gc[1] 0.00985f
C434 PHI_2 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C435 a_23030_n402# EN 0.08752f
C436 VDD a_32570_158# 0.00491f
C437 a_55558_38# gc[10] 0.00972f
C438 a_55214_158# a_55066_158# 0
C439 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_13998_158# 0.01536f
C440 a_45442_n387# a_45198_158# 0.01595f
C441 PHI_1 a_55214_158# 0.01882f
C442 a_11386_158# PHI_1 0.00201f
C443 PHI_1 a_26682_158# 0.00477f
C444 EN a_57882_158# 0.00368f
C445 a_32718_158# VDD 0.55136f
C446 a_7758_158# a_6774_n402# 0.07055f
C447 gc[7] a_35978_n384# 0.00668f
C448 PHI_2 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C449 a_24014_158# PHI_1 0.01882f
C450 PHI_2 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C451 a_13998_158# a_13482_n384# 0.30053f
C452 a_49318_38# VDD 0.32599f
C453 VDD a_26478_158# 0.55136f
C454 a_45050_158# a_45198_158# 0
C455 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_2 0.45413f
C456 a_534_n402# VDD 1.03607f
C457 a_1370_n387# a_1518_158# 0
C458 a_30254_158# a_31734_n402# 0.00268f
C459 a_29270_n402# a_29738_n384# 0.30528f
C460 gc[5] gc[4] 0.01049f
C461 a_13014_n402# PHI_2 0.60119f
C462 a_13850_n387# PHI_2 0
C463 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_35978_n384# 0
C464 EN a_52903_n425# 0.00398f
C465 EN a_51682_n387# 0.00579f
C466 a_42586_n387# a_42218_n384# 0.00194f
C467 PHI_2 a_29738_n384# 0.03321f
C468 a_42978_n387# a_43078_38# 0
C469 PHI_1 a_54230_n402# 0.70141f
C470 a_54698_n384# gc[10] 0.00668f
C471 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_37974_n402# 0
C472 PHI_1 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C473 a_25494_n402# Q[5] 0.00225f
C474 PHI_1 a_26330_158# 0.00164f
C475 EN a_57530_158# 0.00101f
C476 gc[7] a_37974_n402# 0.00985f
C477 a_23030_n402# PHI_1 0.70141f
C478 PHI_2 a_34183_n425# 0
C479 a_48458_n384# VDD 0.4225f
C480 Q[10] gc[10] 0.22358f
C481 PHI_1 a_57882_158# 0.00477f
C482 gc[8] Q[7] 0.17162f
C483 a_29270_n402# a_31734_n402# 0
C484 a_1762_n387# a_1518_158# 0.01595f
C485 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_29738_n384# 0
C486 a_27943_n425# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C487 a_11534_158# PHI_2 0.04895f
C488 gc[4] a_23866_n387# 0
C489 VDD DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42635f
C490 a_34183_n425# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C491 a_14242_n387# PHI_2 0
C492 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_37974_n402# 0.16689f
C493 a_13998_158# VDD 0.55136f
C494 a_54698_n384# a_55558_38# 0.00888f
C495 PHI_2 gc[10] 0.31085f
C496 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD 0.42635f
C497 a_n742_158# a_n946_158# 0.01151f
C498 EN a_55418_158# 0.00368f
C499 a_4310_n402# a_5638_38# 0.02403f
C500 PHI_2 a_31734_n402# 0.60119f
C501 a_1518_158# a_1862_38# 0.57845f
C502 EN D_in 0.13355f
C503 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_21703_n425# 0.0097f
C504 a_30106_158# a_29738_n384# 0.00294f
C505 a_50454_n402# VDD 1.03607f
C506 gc[7] a_36494_158# 0.01329f
C507 PHI_2 a_32570_n387# 0
C508 a_17626_n387# EN 0.0022f
C509 a_17978_158# VDD 0.01506f
C510 PHI_1 a_57530_158# 0.00164f
C511 a_29738_n384# a_30106_n387# 0.00194f
C512 Q[7] PHI_2 0.63578f
C513 a_31734_n402# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C514 Q[3] PHI_2 0.63578f
C515 a_39302_38# a_39162_158# 0.00109f
C516 Q[4] PHI_2 0.63578f
C517 a_29270_n402# a_30254_158# 0.07055f
C518 PHI_2 a_55558_38# 0.03207f
C519 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_31734_n402# 0.16689f
C520 a_24358_38# a_24218_158# 0.00109f
C521 a_42938_158# a_42734_158# 0.01151f
C522 a_30598_38# EN 0.05124f
C523 a_26330_n387# PHI_2 0
C524 a_n1094_158# VDD 0.00491f
C525 Q[8] a_49318_38# 0.00242f
C526 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_36494_158# 0.09501f
C527 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_32570_n387# 0
C528 EN a_55066_158# 0.00101f
C529 a_1370_158# a_1518_158# 0
C530 PHI_2 a_30254_158# 0.04895f
C531 EN PHI_1 0.59089f
C532 a_4310_n402# a_4778_n384# 0.30528f
C533 a_1518_158# a_1002_n384# 0.30053f
C534 gc[2] Q[1] 0.17162f
C535 VDD a_44214_n402# 1.03607f
C536 gc[9] gc[10] 0.01049f
C537 PHI_1 a_55418_158# 0.00534f
C538 a_30458_158# a_30254_158# 0.01151f
C539 Q[1] PHI_2 0.63578f
C540 PHI_2 a_32962_n387# 0
C541 gc[7] a_35510_n402# 0.00985f
C542 D_in PHI_1 0.0221f
C543 a_48974_158# VDD 0.56047f
C544 a_26822_38# a_25962_n384# 0.00888f
C545 gc[8] PHI_2 0.31085f
C546 a_51290_n387# a_50922_n384# 0.00194f
C547 a_17626_158# VDD 0.00491f
C548 a_51682_n387# a_51782_38# 0
C549 Q[9] VDD 0.56326f
C550 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_30254_158# 0.09501f
C551 PHI_2 a_54698_n384# 0.03321f
C552 a_26722_n387# PHI_2 0
C553 a_42586_158# a_42734_158# 0
C554 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_25962_n384# 0
C555 VDD a_45542_38# 0.32599f
C556 a_36698_158# a_36838_38# 0.00109f
C557 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_35510_n402# 0.00116f
C558 Q[8] a_48458_n384# 0.36203f
C559 a_30598_38# PHI_1 0.01314f
C560 PHI_2 Q[10] 0.32019f
C561 PHI_2 a_36838_38# 0.03207f
C562 Q[7] a_37974_n402# 0.00225f
C563 PHI_2 a_29270_n402# 0.02762f
C564 a_4310_n402# a_6774_n402# 0
C565 VDD a_42734_158# 0.56047f
C566 PHI_1 a_55066_158# 0.00201f
C567 gc[2] PHI_2 0.31085f
C568 a_20582_38# EN 0.0522f
C569 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[1] 0.01068f
C570 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_1518_158# 0.00144f
C571 EN a_36346_158# 0.00101f
C572 a_20238_158# VDD 0.55136f
C573 a_30106_158# a_30254_158# 0
C574 EN a_51782_38# 0.0522f
C575 a_n742_158# a_n602_38# 0.00109f
C576 PHI_2 a_36698_158# 0.00411f
C577 a_47990_n402# VDD 1.00028f
C578 a_5498_158# VDD 0.01506f
C579 a_26822_38# a_26478_158# 0.57845f
C580 a_7758_158# a_7962_158# 0.01151f
C581 a_30254_158# a_30106_n387# 0
C582 a_35978_n384# a_36838_38# 0.00888f
C583 a_51290_n387# a_51438_158# 0
C584 a_38958_158# a_39162_158# 0.01151f
C585 gc[8] gc[9] 0.01049f
C586 a_38442_n384# a_38810_158# 0.00294f
C587 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_29270_n402# 0.00116f
C588 a_33062_38# a_31734_n402# 0.02403f
C589 a_30458_158# PHI_2 0.00411f
C590 a_23498_n384# a_23866_158# 0.00294f
C591 VDD a_44682_n384# 0.42245f
C592 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_26478_158# 0.00144f
C593 a_54698_n384# gc[9] 0
C594 a_23030_n402# gc[4] 0.00493f
C595 EN Q[5] 0.513f
C596 PHI_2 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C597 PHI_2 a_35978_n384# 0.03321f
C598 VDD a_41750_n402# 1.00028f
C599 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_2 0.45413f
C600 EN a_5638_38# 0.05124f
C601 gc[8] a_48826_n387# 0
C602 a_19722_n384# EN 0.05124f
C603 a_1722_158# a_1862_38# 0.00109f
C604 PHI_2 a_49218_n387# 0
C605 a_18018_n387# PHI_2 0
C606 EN a_50922_n384# 0.05124f
C607 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[2] 0.23535f
C608 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_534_n402# 0.16689f
C609 a_1518_158# gc[1] 0.01553f
C610 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_2 0.45413f
C611 a_20582_38# PHI_1 0.01261f
C612 a_37974_n402# a_36838_38# 0
C613 a_30254_158# a_30498_n387# 0.01595f
C614 PHI_1 a_36346_158# 0.00201f
C615 a_24358_38# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.2556f
C616 a_51682_n387# a_51438_158# 0.01595f
C617 PHI_1 a_51782_38# 0.01261f
C618 a_38958_158# a_38810_158# 0
C619 a_20238_158# a_20090_n387# 0
C620 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_16790_n402# 0
C621 Q[8] a_44214_n402# 0.00225f
C622 a_32202_n384# a_31734_n402# 0.30528f
C623 PHI_2 gc[9] 0.31085f
C624 a_30106_158# PHI_2 0
C625 Q[1] a_5294_158# 0.01552f
C626 VDD a_45198_158# 0.55136f
C627 a_30598_38# Q[5] 0.00242f
C628 Q[8] a_48974_158# 0.01552f
C629 a_1518_158# VDD 0.55136f
C630 a_32202_n384# a_32570_n387# 0.00194f
C631 a_14342_38# a_14202_158# 0.00109f
C632 PHI_2 a_30106_n387# 0
C633 a_33062_38# a_32962_n387# 0
C634 PHI_2 a_37974_n402# 0.60119f
C635 a_27943_n425# PHI_2 0
C636 Q[5] PHI_1 0.05798f
C637 a_13998_158# gc[3] 0.01553f
C638 EN a_4778_n384# 0.05108f
C639 a_24358_38# VDD 0.32599f
C640 PHI_2 a_48826_n387# 0
C641 EN a_51438_158# 0.11443f
C642 EN a_n946_158# 0.11055f
C643 a_20442_158# PHI_2 0.00422f
C644 Q[8] a_45542_38# 0.25874f
C645 PHI_2 a_51642_158# 0.00422f
C646 a_26330_n387# a_25962_n384# 0.00194f
C647 a_49218_n387# gc[9] 0
C648 PHI_1 a_5638_38# 0.01314f
C649 PHI_1 a_50922_n384# 0.01277f
C650 EN gc[4] 0.44384f
C651 a_37974_n402# a_35978_n384# 0
C652 a_36494_158# a_36838_38# 0.57845f
C653 a_19722_n384# PHI_1 0.01277f
C654 a_23498_n384# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C655 a_n946_158# D_in 0.01538f
C656 Q[2] DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C657 a_32718_158# a_31734_n402# 0.07055f
C658 gc[2] a_5294_158# 0.01329f
C659 VDD a_39162_158# 0.01506f
C660 a_36698_158# a_36494_158# 0.01151f
C661 Q[8] a_47990_n402# 0.16779f
C662 PHI_2 a_5294_158# 0.04895f
C663 PHI_2 a_30498_n387# 0
C664 a_13014_n402# a_13998_158# 0.07055f
C665 a_32718_158# a_32570_n387# 0
C666 PHI_2 a_36494_158# 0.04895f
C667 a_43078_38# a_42938_158# 0.00109f
C668 EN a_10550_n402# 0.08752f
C669 a_13850_n387# a_13998_158# 0
C670 a_33062_38# PHI_2 0.03174f
C671 EN a_6774_n402# 0.08694f
C672 a_17626_n387# gc[4] 0
C673 a_23498_n384# VDD 0.4225f
C674 a_20090_158# PHI_2 0
C675 PHI_2 a_51290_158# 0
C676 gc[6] a_36346_n387# 0
C677 Q[8] a_44682_n384# 0.00101f
C678 a_48826_n387# gc[9] 0
C679 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_51290_n387# 0
C680 a_51642_158# gc[9] 0
C681 PHI_1 a_4778_n384# 0.0533f
C682 a_36494_158# a_35978_n384# 0.30053f
C683 a_35510_n402# a_36838_38# 0.02403f
C684 a_26330_n387# a_26478_158# 0
C685 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_20238_158# 0.01536f
C686 PHI_1 a_51438_158# 0.01804f
C687 a_n946_158# PHI_1 0.01882f
C688 gc[6] VDD 0.26766f
C689 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_33062_38# 0.00242f
C690 gc[4] PHI_1 0.01023f
C691 a_19722_n384# a_20582_38# 0.00888f
C692 a_44214_n402# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.16689f
C693 a_50922_n384# a_51782_38# 0.00888f
C694 VDD a_38810_158# 0.00491f
C695 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_5294_158# 0.09501f
C696 a_13482_n384# a_13850_158# 0.00294f
C697 PHI_2 a_32922_158# 0.00422f
C698 a_32718_158# a_32962_n387# 0.01595f
C699 PHI_2 a_35510_n402# 0.02762f
C700 a_14242_n387# a_13998_158# 0.01595f
C701 a_32202_n384# PHI_2 0.07395f
C702 a_9223_n425# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C703 a_534_n402# Q[1] 0.00225f
C704 PHI_2 a_25962_n384# 0.07395f
C705 PHI_1 a_10550_n402# 0.70141f
C706 Q[8] a_45198_158# 0.11433f
C707 a_58022_38# a_56694_n402# 0.02403f
C708 VDD a_43078_38# 0.32599f
C709 PHI_1 a_6774_n402# 0.01733f
C710 a_35510_n402# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C711 a_36494_158# a_37974_n402# 0.00268f
C712 EN DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C713 a_14202_158# VDD 0.01506f
C714 a_24218_158# gc[5] 0
C715 a_35510_n402# a_35978_n384# 0.30528f
C716 a_26722_n387# a_26478_158# 0.01595f
C717 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_45542_38# 0.00242f
C718 a_32202_n384# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C719 a_1722_158# gc[1] 0
C720 EN a_n602_38# 0.05124f
C721 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_32202_n384# 0.36162f
C722 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_57162_n384# 0
C723 a_7758_158# Q[2] 0.11433f
C724 a_13998_158# Q[3] 0.11433f
C725 a_51438_158# a_51782_38# 0.57845f
C726 a_42734_158# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.09501f
C727 VDD DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42635f
C728 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[4] 0.08575f
C729 PHI_2 a_32570_158# 0
C730 a_n602_38# D_in 0.00242f
C731 a_20582_38# gc[4] 0.01014f
C732 a_42218_n384# a_42586_158# 0.00294f
C733 a_32718_158# PHI_2 0.04011f
C734 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_41750_n402# 0
C735 a_1722_158# VDD 0.01506f
C736 PHI_2 a_49318_38# 0.03207f
C737 gc[8] a_48458_n384# 0
C738 EN DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C739 PHI_2 a_26478_158# 0.04011f
C740 gc[7] a_41750_n402# 0.00493f
C741 gc[1] a_5146_n387# 0
C742 a_534_n402# PHI_2 0.60119f
C743 a_18118_38# EN 0.05124f
C744 a_57162_n384# a_56694_n402# 0.30528f
C745 VDD a_42218_n384# 0.4225f
C746 EN a_48826_158# 0.00101f
C747 EN a_42586_n387# 0.0022f
C748 a_35510_n402# a_37974_n402# 0
C749 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_44682_n384# 0.36162f
C750 a_13850_158# VDD 0.00491f
C751 a_32718_158# DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C752 EN a_n1462_n384# 0.05107f
C753 a_4778_n384# a_5638_38# 0.00888f
C754 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_57678_158# 0.00144f
C755 PHI_1 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C756 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_32718_158# 0.01536f
C757 a_41750_n402# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00116f
C758 a_17774_158# EN 0.11055f
C759 a_51438_158# a_50922_n384# 0.30053f
C760 a_n602_38# PHI_1 0.01314f
C761 Q[9] gc[10] 0.17162f
C762 a_n1462_n384# D_in 0.36155f
C763 Q[6] a_36346_n387# 0
C764 a_49318_38# a_49218_n387# 0
C765 gc[7] a_36738_n387# 0
C766 a_19722_n384# gc[4] 0.00668f
C767 a_5146_158# EN 0.00101f
C768 PHI_2 a_48458_n384# 0.03321f
C769 EN a_46663_n425# 0.00398f
C770 a_17258_n384# EN 0.05108f
C771 a_49318_38# gc[9] 0.00972f
C772 Q[6] VDD 0.56326f
C773 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_58022_38# 0.00242f
C774 a_57678_158# a_56694_n402# 0.07055f
C775 a_17626_n387# a_17774_158# 0
C776 PHI_1 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C777 EN a_42978_n387# 0.00577f
C778 a_18118_38# PHI_1 0.01314f
C779 a_35510_n402# a_36494_158# 0.07055f
C780 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_45198_158# 0.01536f
C781 PHI_2 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C782 a_33062_38# a_32922_158# 0.00109f
C783 Q[9] a_55558_38# 0.00242f
C784 a_6774_n402# a_5638_38# 0
C785 a_13998_158# PHI_2 0.04011f
C786 a_32202_n384# a_33062_38# 0.00888f
C787 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_1518_158# 0.01536f
C788 a_57882_158# a_58022_38# 0.00109f
C789 PHI_1 a_48826_158# 0.00201f
C790 a_16790_n402# EN 0.08752f
C791 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C792 a_n1462_n384# PHI_1 0.0533f
C793 gc[8] a_44214_n402# 0.00985f
C794 a_17626_n387# a_17258_n384# 0.00194f
C795 a_7758_158# VDD 0.55136f
C796 Q[7] a_42734_158# 0.01552f
C797 a_17774_158# PHI_1 0.01882f
C798 gc[7] a_39162_158# 0
C799 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_13482_n384# 0
C800 a_7242_n384# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C801 PHI_2 a_50454_n402# 0.60119f
C802 EN a_45050_n387# 0.0022f
C803 a_7610_n387# a_7758_158# 0
C804 a_20238_158# Q[4] 0.11433f
C805 a_17978_158# PHI_2 0.00411f
C806 a_48458_n384# gc[9] 0.00668f
C807 a_19254_n402# EN 0.08694f
C808 EN a_7962_158# 0.00368f
C809 gc[5] DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.23535f
C810 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_57162_n384# 0.36162f
C811 a_5146_158# PHI_1 0.00201f
C812 a_11386_n387# Q[2] 0
C813 a_17258_n384# PHI_1 0.0533f
C814 a_2983_n425# EN 0.00398f
C815 EN a_45402_158# 0.00368f
C816 gc[8] a_45542_38# 0.01014f
C817 a_n1094_158# PHI_2 0
C818 a_6774_n402# a_4778_n384# 0
C819 Q[9] a_54698_n384# 0.36203f
C820 a_24218_158# a_24014_158# 0.01151f
C821 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gc[9] 0.33472f
C822 a_32718_158# a_33062_38# 0.57845f
C823 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_51782_38# 0.00242f
C824 gc[8] a_42734_158# 0.01329f
C825 PHI_2 a_44214_n402# 0.60119f
C826 gc[6] gc[7] 0.01049f
C827 a_48458_n384# a_48826_n387# 0.00194f
C828 Q[7] a_41750_n402# 0.16779f
C829 a_16790_n402# PHI_1 0.70141f
C830 gc[5] VDD 0.26766f
C831 a_7758_158# a_8102_38# 0.57845f
C832 PHI_2 a_48974_158# 0.04895f
C833 gc[8] a_47990_n402# 0.00493f
C834 EN a_45442_n387# 0.00579f
C835 a_8002_n387# a_7758_158# 0.01595f
C836 EN a_58022_38# 0.0522f
C837 a_17626_158# PHI_2 0
C838 a_50454_n402# gc[9] 0.00985f
C839 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_57678_158# 0.01536f
C840 Q[9] PHI_2 0.63578f
C841 EN a_45050_158# 0.00101f
C842 a_32718_158# a_32922_158# 0.01151f
C843 a_1370_n387# EN 0.0022f
C844 a_19254_n402# PHI_1 0.01733f
C845 a_32202_n384# a_32570_158# 0.00294f
C846 PHI_1 a_7962_158# 0.00477f
C847 gc[8] a_44682_n384# 0.00668f
C848 PHI_2 a_45542_38# 0.03174f
C849 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD 0.42635f
C850 a_23866_158# a_24014_158# 0
C851 a_57530_158# a_57162_n384# 0.00294f
C852 a_32718_158# a_32202_n384# 0.30053f
C853 a_57882_158# a_57678_158# 0.01151f
C854 PHI_1 a_45402_158# 0.00477f
C855 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_50922_n384# 0.36162f
C856 a_14202_158# gc[3] 0
C857 PHI_2 a_42734_158# 0.04895f
C858 gc[8] a_41750_n402# 0.00985f
C859 a_5498_158# gc[2] 0
C860 a_26478_158# a_25962_n384# 0.30053f
C861 a_48974_158# a_49218_n387# 0.01595f
C862 a_n742_158# gc[1] 0
C863 gc[6] a_29738_n384# 0.00668f
C864 a_43078_38# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.2556f
C865 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_4310_n402# 0
C866 a_n946_158# a_n602_38# 0.57845f
C867 a_24358_38# Q[4] 0.00242f
C868 a_20238_158# PHI_2 0.04011f
C869 EN a_57162_n384# 0.05124f
C870 a_7758_158# a_7242_n384# 0.30053f
C871 PHI_2 a_47990_n402# 0.02762f
C872 a_5498_158# PHI_2 0.00411f
C873 EN a_49178_158# 0.00368f
C874 a_7610_158# VDD 0.00491f
C875 a_48974_158# gc[9] 0.01329f
C876 a_20482_n387# EN 0.00579f
C877 VDD DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.4236f
C878 gc[6] a_34183_n425# 0.00113f
C879 PHI_1 a_58022_38# 0.01261f
C880 a_25494_n402# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.16689f
C881 a_1762_n387# EN 0.00579f
C882 a_n742_158# VDD 0.01506f
C883 a_32718_158# a_32570_158# 0
C884 a_1518_158# Q[1] 0.11433f
C885 Q[9] gc[9] 0.22418f
C886 gc[7] a_42218_n384# 0
C887 PHI_2 a_44682_n384# 0.07395f
C888 gc[8] a_45198_158# 0.01553f
C889 EN a_39302_38# 0.0522f
C890 a_57530_158# a_57678_158# 0
C891 PHI_1 a_45050_158# 0.00164f
C892 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_51438_158# 0.01536f
C893 a_20582_38# a_19254_n402# 0.02403f
C894 PHI_2 a_41750_n402# 0.02762f
C895 a_48974_158# a_48826_n387# 0
C896 VDD a_56694_n402# 1.03607f
C897 a_1862_38# EN 0.0522f
C898 gc[6] a_31734_n402# 0.00985f
C899 a_18118_38# gc[4] 0.00972f
C900 a_42218_n384# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C901 a_n946_158# a_n1462_n384# 0.30053f
C902 a_36738_n387# a_36838_38# 0
C903 gc[1] a_4310_n402# 0.00493f
C904 a_23498_n384# Q[4] 0.36203f
C905 EN a_57678_158# 0.11443f
C906 a_25494_n402# VDD 1.03607f
C907 a_24218_158# EN 0.00368f
C908 a_47990_n402# gc[9] 0.00985f
C909 a_59143_n425# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C910 gc[6] a_32570_n387# 0
C911 EN a_n1930_n402# 0.08666f
C912 PHI_1 a_57162_n384# 0.01277f
C913 PHI_1 a_49178_158# 0.00534f
C914 Q[6] gc[7] 0.17162f
C915 EN a_38810_n387# 0.0022f
C916 a_24014_158# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.09501f
C917 a_17774_158# gc[4] 0.01329f
C918 PHI_2 a_45198_158# 0.04011f
C919 EN a_38442_n384# 0.05124f
C920 a_5146_158# a_4778_n384# 0.00294f
C921 PHI_2 a_36738_n387# 0
C922 VDD a_4310_n402# 1.00028f
C923 a_1518_158# PHI_2 0.04011f
C924 D_in a_n1930_n402# 0.15891f
C925 a_19722_n384# a_19254_n402# 0.30528f
C926 a_48458_n384# a_49318_38# 0.00888f
C927 PHI_1 a_39302_38# 0.01261f
C928 a_20442_158# a_20238_158# 0.01151f
C929 a_1370_158# EN 0.00101f
C930 VDD a_55214_158# 0.56047f
C931 a_24358_38# PHI_2 0.03207f
C932 Q[6] DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C933 a_1002_n384# EN 0.05124f
C934 VDD a_26682_158# 0.01506f
C935 a_17258_n384# gc[4] 0.00668f
C936 gc[6] a_30254_158# 0.01329f
C937 a_11386_158# VDD 0.00491f
C938 a_24014_158# VDD 0.56047f
C939 Q[7] a_43078_38# 0.00242f
C940 a_1862_38# PHI_1 0.01261f
C941 a_14342_38# EN 0.0522f
C942 a_23866_158# EN 0.00101f
C943 gc[6] a_32962_n387# 0
C944 PHI_1 a_57678_158# 0.01804f
C945 EN a_39202_n387# 0.00579f
C946 a_7242_n384# a_7610_158# 0.00294f
C947 a_23030_n402# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00116f
C948 a_16790_n402# gc[4] 0.00985f
C949 a_24218_158# PHI_1 0.00534f
C950 EN a_38958_158# 0.11443f
C951 EN Q[2] 0.513f
C952 PHI_2 a_39162_158# 0.00422f
C953 PHI_1 a_n1930_n402# 0.70141f
C954 a_5498_158# a_5294_158# 0.01151f
C955 a_20482_n387# a_20582_38# 0
C956 PHI_1 a_38442_n384# 0.01277f
C957 a_50454_n402# a_49318_38# 0
C958 a_20090_158# a_20238_158# 0
C959 Q[6] a_34183_n425# 0.00241f
C960 VDD DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C961 VDD a_54230_n402# 1.00028f
C962 a_23498_n384# PHI_2 0.03321f
C963 gc[6] a_29270_n402# 0.00985f
C964 gc[5] a_26822_38# 0.01014f
C965 a_19254_n402# gc[4] 0.00985f
C966 VDD a_26330_158# 0.00491f
C967 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q EN 0.20415f
C968 a_1370_158# PHI_1 0.00164f
C969 gc[8] a_43078_38# 0.00972f
C970 a_23030_n402# VDD 1.00028f
C971 a_1002_n384# PHI_1 0.01277f
C972 Q[7] a_42218_n384# 0.36203f
C973 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN 0.65271f
C974 a_13482_n384# EN 0.05124f
C975 VDD a_57882_158# 0.01506f
C976 gc[5] DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.33472f
C977 a_n1462_n384# a_n602_38# 0.00888f
C978 gc[6] PHI_2 0.31085f
C979 EN a_42938_158# 0.00368f
C980 a_14342_38# PHI_1 0.01261f
C981 a_23866_158# PHI_1 0.00201f
C982 PHI_2 a_38810_158# 0
C983 Q[6] a_31734_n402# 0.00225f
C984 a_30458_158# gc[6] 0
C985 a_15463_n425# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C986 a_50454_n402# a_48458_n384# 0
C987 PHI_1 a_38958_158# 0.01804f
C988 a_48974_158# a_49318_38# 0.57845f
C989 Q[2] PHI_1 0.05798f
C990 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gc[3] 0.33472f
C991 gc[6] DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.33472f
C992 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_46663_n425# 0.0097f
C993 gc[6] a_35978_n384# 0
C994 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[6] 0.23535f
C995 a_9223_n425# EN 0.00398f
C996 a_36738_n387# a_36494_158# 0.01595f
C997 EN DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C998 gc[8] a_42218_n384# 0.00668f
C999 PHI_2 a_43078_38# 0.03207f
C1000 a_n1094_n387# EN 0.0022f
C1001 a_50454_n402# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1002 a_14202_158# PHI_2 0.00422f
C1003 a_18118_38# a_17774_158# 0.57845f
C1004 EN gc[1] 0.44384f
C1005 gc[5] a_29738_n384# 0
C1006 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_1 0.01369f
C1007 VDD a_57530_158# 0.00491f
C1008 Q[1] a_5146_n387# 0
C1009 gc[2] DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.33472f
C1010 EN a_42586_158# 0.00101f
C1011 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C1012 EN a_36346_n387# 0.0022f
C1013 a_13482_n384# PHI_1 0.01277f
C1014 a_n1094_n387# D_in 0
C1015 a_11018_n384# a_11386_n387# 0.00194f
C1016 a_13014_n402# DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1017 PHI_2 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C1018 a_11878_38# a_11778_n387# 0
C1019 gc[1] D_in 0.17162f
C1020 PHI_1 a_42938_158# 0.00534f
C1021 a_17258_n384# a_18118_38# 0.00888f
C1022 a_48974_158# a_48458_n384# 0.30053f
C1023 a_47990_n402# a_49318_38# 0.02403f
C1024 EN VDD 3.51464f
C1025 a_11386_n387# gc[3] 0
C1026 a_1722_158# PHI_2 0.00422f
C1027 gc[6] a_30106_n387# 0
C1028 a_57530_n387# DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C1029 a_7610_n387# EN 0.0022f
C1030 VDD a_55418_158# 0.01506f
C1031 a_20482_n387# gc[4] 0
C1032 EN a_21703_n425# 0.00398f
C1033 PHI_2 a_42218_n384# 0.03321f
C1034 a_25494_n402# a_26822_38# 0.02403f
C1035 D_in VDD 0.18307f
C1036 EN a_40423_n425# 0.00398f
C1037 a_n702_n387# EN 0.00577f
C1038 a_18118_38# a_16790_n402# 0.02403f
C1039 a_17258_n384# a_17774_158# 0.30053f
C1040 a_13850_158# PHI_2 0
C1041 PHI_1 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C1042 gc[2] a_5146_n387# 0
C1043 Q[9] DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1044 gc[1] PHI_1 0.01023f
C1045 a_25494_n402# DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1046 PHI_2 a_5146_n387# 0
C1047 Q[6] a_36838_38# 0.00242f
C1048 PHI_1 a_42586_158# 0.00201f
C1049 a_30598_38# VDD 0.32599f
C1050 a_16790_n402# a_17774_158# 0.07055f
C1051 a_19254_n402# a_18118_38# 0
C1052 a_47990_n402# a_48458_n384# 0.30528f
C1053 a_48974_158# a_50454_n402# 0.00268f
C1054 EN a_59143_n425# 0.00398f
C1055 a_11778_n387# gc[3] 0
C1056 gc[5] Q[4] 0.17162f
C1057 a_n946_158# a_n1930_n402# 0.07055f
C1058 gc[6] a_30498_n387# 0
C1059 a_8102_38# EN 0.0522f
C1060 a_26330_n387# gc[5] 0
C1061 a_8002_n387# EN 0.00579f
C1062 Q[9] a_50454_n402# 0.00225f
C1063 a_26822_38# a_26682_158# 0.00109f
C1064 a_33062_38# gc[6] 0.01014f
C1065 a_11018_n384# a_11386_158# 0.00294f
C1066 VDD a_55066_158# 0.00491f
C1067 PHI_1 VDD 9.88453f
C1068 EN a_20090_n387# 0.0022f
C1069 Q[6] PHI_2 0.63578f
C1070 a_19254_n402# a_17774_158# 0.00268f
C1071 a_17258_n384# a_16790_n402# 0.30528f
C1072 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_20238_158# 0.00144f
C1073 gc[2] a_5538_n387# 0
C1074 a_1518_158# a_534_n402# 0.07055f
C1075 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[3] 0.08575f
C1076 a_7758_158# gc[2] 0.01553f
C1077 Q[6] DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1078 PHI_2 a_5538_n387# 0
C1079 Q[6] a_35978_n384# 0.36203f
C1080 a_11534_158# a_11386_n387# 0
C1081 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gc[10] 0.33472f
C1082 a_7758_158# PHI_2 0.04011f
C1083 a_19254_n402# a_17258_n384# 0
C1084 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[6] 0.01102f
C1085 EN a_57530_n387# 0.0022f
C1086 a_47990_n402# a_50454_n402# 0
C1087 gc[6] a_32922_158# 0
C1088 gc[6] a_35510_n402# 0.00493f
C1089 Q[4] a_23866_n387# 0
C1090 a_44214_n402# a_45542_38# 0.02403f
C1091 a_7242_n384# EN 0.05124f
C1092 a_26722_n387# gc[5] 0
C1093 a_32202_n384# gc[6] 0.00668f
C1094 a_11738_158# EN 0.00368f
C1095 Q[5] DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01102f
C1096 a_19254_n402# a_16790_n402# 0
C1097 a_8102_38# PHI_1 0.01261f
C1098 a_56694_n402# gc[10] 0.00985f
C1099 a_42734_158# a_44214_n402# 0.00268f
C1100 gc[5] a_29270_n402# 0.00493f
C1101 VDD a_36346_158# 0.00491f
C1102 VDD a_51782_38# 0.32599f
C1103 EN Q[8] 0.513f
C1104 a_20582_38# VDD 0.32599f
C1105 a_55066_n387# gc[10] 0
C1106 a_11534_158# a_11778_n387# 0.01595f
C1107 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_7758_158# 0.01536f
C1108 gc[5] PHI_2 0.31085f
C1109 a_47990_n402# a_48974_158# 0.07055f
C1110 EN a_57922_n387# 0.00579f
C1111 a_11878_38# EN 0.05124f
C1112 Q[2] a_10550_n402# 0.16779f
C1113 Q[5] VDD 0.56326f
C1114 a_56694_n402# a_55558_38# 0
C1115 a_44214_n402# a_44682_n384# 0.30528f
C1116 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q EN 0.20415f
C1117 a_5146_n387# a_5294_158# 0
C1118 Q[2] a_6774_n402# 0.00225f
C1119 a_32718_158# gc[6] 0.01553f
C1120 a_11534_158# a_11386_158# 0
C1121 a_7242_n384# PHI_1 0.01277f
C1122 a_n602_38# a_n1930_n402# 0.02403f
C1123 a_55214_158# gc[10] 0.01329f
C1124 VDD a_5638_38# 0.32599f
C1125 a_41750_n402# a_44214_n402# 0
C1126 a_19722_n384# VDD 0.42245f
C1127 a_11738_158# PHI_1 0.00534f
C1128 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_10550_n402# 0.00116f
C1129 VDD a_50922_n384# 0.42245f
C1130 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C1131 Q[8] PHI_1 0.05798f
C1132 a_55458_n387# gc[10] 0
C1133 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q[10] 0.08537f
C1134 Q[6] a_36494_158# 0.01552f
C1135 a_44682_n384# a_45542_38# 0.00888f
C1136 a_n1094_n387# a_n946_158# 0
C1137 a_33062_38# Q[6] 0.25874f
C1138 gc[1] a_4778_n384# 0
C1139 EN DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C1140 PHI_2 a_23866_n387# 0
C1141 a_n946_158# gc[1] 0.01329f
C1142 a_11018_n384# EN 0.05108f
C1143 EN a_26822_38# 0.0522f
C1144 EN gc[7] 0.44384f
C1145 a_15463_n425# EN 0.00398f
C1146 a_56694_n402# a_54698_n384# 0
C1147 a_55214_158# a_55558_38# 0.57845f
C1148 a_44214_n402# a_45198_158# 0.07055f
C1149 a_7610_158# PHI_2 0
C1150 a_5538_n387# a_5294_158# 0.01595f
C1151 a_11878_38# PHI_1 0.01314f
C1152 gc[3] EN 0.44384f
C1153 a_24014_158# Q[4] 0.01552f
C1154 PHI_2 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C1155 a_11386_n387# gc[2] 0
C1156 EN DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C1157 Q[1] a_4310_n402# 0.16779f
C1158 a_n1462_n384# a_n1930_n402# 0.30528f
C1159 a_56694_n402# Q[10] 0.00225f
C1160 VDD a_4778_n384# 0.4225f
C1161 gc[5] a_30106_n387# 0
C1162 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_1 0.01369f
C1163 a_54230_n402# gc[10] 0.00985f
C1164 a_41750_n402# a_42734_158# 0.07055f
C1165 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[10] 0.23535f
C1166 a_n742_158# PHI_2 0.00411f
C1167 a_55066_n387# a_54698_n384# 0.00194f
C1168 a_n946_158# VDD 0.56047f
C1169 VDD a_51438_158# 0.55136f
C1170 a_55458_n387# a_55558_38# 0
C1171 a_11386_n387# PHI_2 0
C1172 a_27943_n425# gc[5] 0.00113f
C1173 EN DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C1174 EN DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C1175 gc[4] VDD 0.26766f
C1176 Q[6] a_35510_n402# 0.16779f
C1177 a_57882_158# gc[10] 0
C1178 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q EN 0.20415f
C1179 a_19722_n384# a_20090_n387# 0.00194f
C1180 a_32202_n384# Q[6] 0.00101f
C1181 a_45198_158# a_45542_38# 0.57845f
C1182 a_n702_n387# a_n946_158# 0.01595f
C1183 a_17626_n387# gc[3] 0
C1184 PHI_2 a_56694_n402# 0.60119f
C1185 PHI_2 a_24258_n387# 0
C1186 a_13014_n402# EN 0.08694f
C1187 gc[4] a_21703_n425# 0.00113f
C1188 a_25494_n402# PHI_2 0.60119f
C1189 a_54230_n402# a_55558_38# 0.02403f
C1190 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q D_in 0.01068f
C1191 a_55214_158# a_54698_n384# 0.30053f
C1192 a_13850_n387# EN 0.0022f
C1193 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_55558_38# 0.2556f
C1194 PHI_1 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C1195 VDD a_10550_n402# 1.00028f
C1196 a_11018_n384# PHI_1 0.0533f
C1197 a_23030_n402# Q[4] 0.16779f
C1198 PHI_1 a_26822_38# 0.01261f
C1199 PHI_2 a_55066_n387# 0
C1200 EN a_29738_n384# 0.05108f
C1201 gc[7] PHI_1 0.01023f
C1202 gc[2] a_4310_n402# 0.00985f
C1203 VDD a_6774_n402# 1.03607f
C1204 gc[3] PHI_1 0.01023f
C1205 a_11778_n387# PHI_2 0
C1206 PHI_1 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C1207 PHI_2 a_4310_n402# 0.02762f
C1208 EN a_34183_n425# 0.00398f
C1209 a_13998_158# a_14202_158# 0.01151f
C1210 a_20582_38# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00242f
C1211 a_57162_n384# a_58022_38# 0.00888f
C1212 a_45198_158# a_44682_n384# 0.30053f
C1213 a_32718_158# Q[6] 0.11433f
C1214 PHI_1 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C1215 PHI_2 a_55214_158# 0.04895f
C1216 PHI_1 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C1217 a_11534_158# EN 0.11055f
C1218 PHI_2 a_26682_158# 0.00422f
C1219 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_1 0.01369f
C1220 a_11386_158# PHI_2 0
C1221 gc[4] a_20090_n387# 0
C1222 a_14242_n387# EN 0.00579f
C1223 a_54230_n402# a_54698_n384# 0.30528f
C1224 a_24014_158# PHI_2 0.04895f
C1225 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_54698_n384# 0
C1226 EN gc[10] 0.4397f
C1227 a_13014_n402# PHI_1 0.01733f
C1228 a_n602_38# gc[1] 0.00972f
C1229 PHI_2 a_55458_n387# 0
C1230 a_30598_38# a_29738_n384# 0.00888f
C1231 EN a_31734_n402# 0.08694f
C1232 a_55066_n387# gc[9] 0
C1233 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[10] 0.01102f
C1234 a_55418_158# gc[10] 0
C1235 PHI_1 a_29738_n384# 0.0533f
C1236 a_8102_38# a_6774_n402# 0.02403f
C1237 EN a_32570_n387# 0.0022f
C1238 a_13998_158# a_13850_158# 0
C1239 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_4310_n402# 0.00116f
C1240 a_19722_n384# DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.36162f
C1241 gc[5] a_25962_n384# 0.00668f
C1242 a_43078_38# a_44214_n402# 0
C1243 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD 0.42635f
C1244 a_57678_158# a_58022_38# 0.57845f
C1245 EN Q[7] 0.513f
C1246 a_n602_38# VDD 0.32599f
C1247 EN Q[4] 0.513f
C1248 PHI_2 a_54230_n402# 0.02762f
C1249 Q[3] EN 0.513f
C1250 PHI_2 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C1251 EN a_55558_38# 0.05124f
C1252 a_26330_n387# EN 0.0022f
C1253 PHI_2 a_26330_158# 0
C1254 PHI_2 a_51290_n387# 0
C1255 Q[5] a_26822_38# 0.25874f
C1256 a_23030_n402# PHI_2 0.02762f
C1257 a_n702_n387# a_n602_38# 0
C1258 a_n1094_n387# a_n1462_n384# 0.00194f
C1259 a_11534_158# PHI_1 0.01882f
C1260 a_55558_38# a_55418_158# 0.00109f
C1261 a_n1462_n384# gc[1] 0.00668f
C1262 a_30598_38# a_31734_n402# 0
C1263 PHI_2 a_57882_158# 0.00422f
C1264 EN a_30254_158# 0.11055f
C1265 Q[5] DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1266 VDD DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C1267 PHI_1 gc[10] 0.00846f
C1268 a_18118_38# VDD 0.32599f
C1269 EN Q[1] 0.513f
C1270 a_17626_n387# Q[3] 0
C1271 PHI_1 a_31734_n402# 0.01733f
C1272 a_7242_n384# a_6774_n402# 0.30528f
C1273 a_48826_158# VDD 0.00491f
C1274 EN a_32962_n387# 0.00579f
C1275 gc[5] a_26478_158# 0.01553f
C1276 a_43078_38# a_42734_158# 0.57845f
C1277 a_42218_n384# a_44214_n402# 0
C1278 a_57678_158# a_57162_n384# 0.30053f
C1279 a_n1462_n384# VDD 0.4225f
C1280 EN gc[8] 0.44384f
C1281 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q gc[4] 0.23535f
C1282 a_1762_n387# a_1862_38# 0
C1283 a_1370_n387# a_1002_n384# 0.00194f
C1284 EN a_54698_n384# 0.05108f
C1285 PHI_2 a_52903_n425# 0
C1286 a_4310_n402# a_5294_158# 0.07055f
C1287 a_26722_n387# EN 0.00579f
C1288 a_17774_158# VDD 0.56047f
C1289 PHI_2 a_51682_n387# 0
C1290 Q[7] PHI_1 0.05798f
C1291 a_54230_n402# gc[9] 0.00493f
C1292 Q[4] PHI_1 0.05798f
C1293 Q[3] PHI_1 0.05798f
C1294 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_2983_n425# 0.0097f
C1295 a_51290_n387# gc[9] 0
C1296 PHI_1 a_55558_38# 0.01314f
C1297 EN Q[10] 0.38669f
C1298 PHI_2 a_57530_158# 0
C1299 a_11878_38# a_10550_n402# 0.02403f
C1300 EN a_36838_38# 0.05124f
C1301 a_30598_38# a_30254_158# 0.57845f
C1302 EN a_29270_n402# 0.08752f
C1303 a_5146_158# VDD 0.00491f
C1304 Q[5] a_29738_n384# 0.36203f
C1305 a_17258_n384# VDD 0.4225f
C1306 PHI_1 a_30254_158# 0.01882f
C1307 gc[2] EN 0.44384f
C1308 a_38442_n384# a_39302_38# 0.00888f
C1309 EN a_36698_158# 0.00368f
C1310 a_23498_n384# a_24358_38# 0.00888f
C1311 a_43078_38# a_41750_n402# 0.02403f
C1312 a_42218_n384# a_42734_158# 0.30053f
C1313 EN PHI_2 1.35356f
C1314 Q[1] PHI_1 0.05798f
C1315 a_25494_n402# a_25962_n384# 0.30528f
C1316 a_16790_n402# VDD 1.00028f
C1317 PHI_2 a_55418_158# 0.00411f
C1318 gc[3] gc[4] 0.01049f
C1319 gc[8] PHI_1 0.01023f
C1320 a_30458_158# EN 0.00368f
C1321 a_52903_n425# gc[9] 0.00113f
C1322 a_51682_n387# gc[9] 0
C1323 D_in PHI_2 0.34149f
C1324 a_2983_n425# gc[1] 0.00113f
C1325 PHI_1 a_54698_n384# 0.0533f
C1326 Q[8] DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1327 EN DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C1328 a_11018_n384# a_10550_n402# 0.30528f
C1329 a_54698_n384# a_55066_158# 0.00294f
C1330 EN a_35978_n384# 0.05108f
C1331 a_30598_38# a_29270_n402# 0.02403f
C1332 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_n946_158# 0.09501f
C1333 a_1002_n384# a_1862_38# 0.00888f
C1334 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q EN 0.20415f
C1335 a_20582_38# Q[4] 0.25874f
C1336 a_17626_n387# PHI_2 0
C1337 a_19254_n402# VDD 1.03607f
C1338 PHI_1 Q[10] 0.03331f
C1339 PHI_1 a_36838_38# 0.01314f
C1340 a_39302_38# a_39202_n387# 0
C1341 a_38442_n384# a_38810_n387# 0.00194f
C1342 gc[3] a_10550_n402# 0.00985f
C1343 VDD a_7962_158# 0.01506f
C1344 PHI_1 a_29270_n402# 0.70141f
C1345 a_38958_158# a_39302_38# 0.57845f
C1346 EN a_49218_n387# 0.00577f
C1347 a_18018_n387# EN 0.00577f
C1348 a_42218_n384# a_41750_n402# 0.30528f
C1349 a_45402_158# VDD 0.01506f
C1350 a_30598_38# PHI_2 0.03207f
C1351 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_13998_158# 0.00144f
C1352 gc[2] PHI_1 0.01023f
C1353 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q EN 0.20415f
C1354 a_25494_n402# a_26478_158# 0.07055f
C1355 PHI_1 a_36698_158# 0.00534f
C1356 EN gc[9] 0.44384f
C1357 Q[8] DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C1358 PHI_2 a_55066_158# 0
C1359 a_30598_38# a_30458_158# 0.00109f
C1360 PHI_2 PHI_1 24.2698f
C1361 a_30106_158# EN 0.00101f
C1362 a_1370_n387# gc[1] 0
C1363 a_13014_n402# a_10550_n402# 0
C1364 EN a_30106_n387# 0.0022f
C1365 EN a_37974_n402# 0.08694f
C1366 a_30458_158# PHI_1 0.00534f
C1367 a_1722_158# a_1518_158# 0.01151f
C1368 a_1370_158# a_1002_n384# 0.00294f
C1369 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_30598_38# 0.2556f
C1370 VDD a_58022_38# 0.32599f
C1371 a_19722_n384# Q[4] 0.00101f
C1372 Q[5] a_30254_158# 0.01552f
C1373 a_27943_n425# EN 0.00398f
C1374 a_38958_158# a_38810_n387# 0
C1375 PHI_1 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C1376 PHI_1 a_35978_n384# 0.0533f
C1377 EN a_48826_n387# 0.0022f
C1378 EN a_51642_158# 0.00368f
C1379 a_20442_158# EN 0.00368f
C1380 a_38958_158# a_38442_n384# 0.30053f
C1381 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_1 0.01369f
C1382 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_18118_38# 0.2556f
C1383 a_45050_158# VDD 0.00491f
C1384 a_26330_158# a_25962_n384# 0.00294f
C1385 a_8102_38# a_7962_158# 0.00109f
C1386 a_26682_158# a_26478_158# 0.01151f
C1387 Q[8] a_46663_n425# 0.00241f
C1388 Q[1] a_5638_38# 0.00242f
C1389 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q PHI_1 0.01369f
C1390 PHI_1 gc[9] 0.01023f
C1391 a_1762_n387# gc[1] 0
C1392 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_17774_158# 0.09501f
C1393 EN a_5294_158# 0.11055f
C1394 EN a_30498_n387# 0.00577f
C1395 a_30106_158# PHI_1 0.00201f
C1396 a_11534_158# a_10550_n402# 0.07055f
C1397 PHI_2 a_36346_158# 0
C1398 PHI_2 a_51782_38# 0.03174f
C1399 a_20582_38# PHI_2 0.03174f
C1400 EN a_36494_158# 0.11055f
C1401 a_33062_38# EN 0.0522f
C1402 VDD a_57162_n384# 0.42245f
C1403 Q[5] a_29270_n402# 0.16779f
C1404 VDD a_49178_158# 0.01506f
C1405 a_38958_158# a_39202_n387# 0.01595f
C1406 PHI_1 a_37974_n402# 0.01733f
C1407 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_n602_38# 0.2556f
C1408 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_1002_n384# 0
C1409 EN a_51290_158# 0.00101f
C1410 a_20090_158# EN 0.00101f
C1411 Q[4] gc[4] 0.22418f
C1412 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_17258_n384# 0
C1413 Q[3] gc[4] 0.17162f
C1414 a_1862_38# gc[1] 0.01014f
C1415 a_26330_158# a_26478_158# 0
C1416 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_14342_38# 0.00242f
C1417 a_35978_n384# a_36346_158# 0.00294f
C1418 VDD a_39302_38# 0.32599f
C1419 PHI_1 a_51642_158# 0.00477f
C1420 a_20442_158# PHI_1 0.00477f
C1421 Q[5] PHI_2 0.63578f
C1422 gc[7] a_42586_n387# 0
C1423 a_13482_n384# a_14342_38# 0.00888f
C1424 gc[2] a_5638_38# 0.00972f
C1425 Q[1] a_4778_n384# 0.36203f
C1426 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[2] 0.01068f
C1427 gc[1] a_n1930_n402# 0.00985f
C1428 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_16790_n402# 0.00116f
C1429 a_1862_38# VDD 0.32599f
C1430 PHI_2 a_5638_38# 0.03207f
C1431 a_30598_38# a_30498_n387# 0
C1432 EN a_32922_158# 0.00368f
C1433 a_19722_n384# PHI_2 0.07395f
C1434 EN a_35510_n402# 0.08752f
C1435 PHI_2 a_50922_n384# 0.07395f
C1436 VDD a_57678_158# 0.55136f
C1437 a_32202_n384# EN 0.05124f
C1438 a_51782_38# gc[9] 0.01014f
C1439 PHI_1 a_5294_158# 0.01882f
C1440 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q Q[5] 0.01068f
C1441 PHI_1 a_36494_158# 0.01882f
C1442 EN a_25962_n384# 0.05124f
C1443 a_24218_158# VDD 0.01506f
C1444 VDD a_n1930_n402# 0.99746f
C1445 a_33062_38# PHI_1 0.01261f
C1446 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_n1462_n384# 0
C1447 a_1002_n384# gc[1] 0.00668f
C1448 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_19254_n402# 0.16689f
C1449 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_13482_n384# 0.36162f
C1450 a_17258_n384# gc[3] 0
C1451 a_20090_158# PHI_1 0.00164f
C1452 VDD a_38442_n384# 0.42245f
C1453 PHI_1 a_51290_158# 0.00164f
C1454 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_54230_n402# 0
C1455 gc[2] a_4778_n384# 0.00668f
C1456 a_42218_n384# a_43078_38# 0.00888f
C1457 a_20582_38# a_20442_158# 0.00109f
C1458 a_9223_n425# Q[2] 0.00241f
C1459 a_51782_38# a_51642_158# 0.00109f
C1460 a_1370_158# VDD 0.00491f
C1461 a_1002_n384# VDD 0.42245f
C1462 PHI_2 a_4778_n384# 0.03321f
C1463 Q[9] a_55066_n387# 0
C1464 EN a_32570_158# 0.00101f
C1465 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_5638_38# 0.2556f
C1466 Q[6] gc[6] 0.22418f
C1467 a_16790_n402# gc[3] 0.00493f
C1468 Q[5] a_30106_n387# 0
C1469 a_n946_158# PHI_2 0.04895f
C1470 PHI_2 a_51438_158# 0.04011f
C1471 a_57922_n387# a_58022_38# 0
C1472 a_57530_n387# a_57162_n384# 0.00194f
C1473 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_23030_n402# 0
C1474 a_32718_158# EN 0.11443f
C1475 PHI_1 a_32922_158# 0.00477f
C1476 EN a_49318_38# 0.05124f
C1477 a_50922_n384# gc[9] 0.00668f
C1478 a_27943_n425# Q[5] 0.00241f
C1479 a_24358_38# gc[5] 0.00972f
C1480 a_14342_38# VDD 0.32599f
C1481 PHI_1 a_35510_n402# 0.70141f
C1482 gc[4] PHI_2 0.31085f
C1483 a_23866_158# VDD 0.00491f
C1484 EN a_26478_158# 0.11443f
C1485 EN a_534_n402# 0.08694f
C1486 a_32202_n384# PHI_1 0.01277f
C1487 PHI_1 a_25962_n384# 0.01277f
C1488 a_36494_158# a_36346_158# 0
C1489 gc[2] a_10550_n402# 0.00493f
C1490 VDD a_38958_158# 0.55136f
C1491 Q[9] a_55214_158# 0.01552f
C1492 Q[2] VDD 0.56326f
C1493 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gc[1] 0.33472f
C1494 PHI_2 a_10550_n402# 0.02762f
C1495 gc[2] a_6774_n402# 0.00985f
C1496 a_52903_n425# DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C1497 a_45050_n387# DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C1498 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_4778_n384# 0
C1499 PHI_2 a_6774_n402# 0.60119f
C1500 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD 0.34237f
C1501 a_18018_n387# gc[4] 0
C1502 a_51438_158# gc[9] 0.01553f
C1503 a_57530_n387# a_57678_158# 0
C1504 a_18118_38# Q[3] 0.00242f
C1505 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD 0.42635f
C1506 EN a_48458_n384# 0.05108f
C1507 a_23498_n384# gc[5] 0.00668f
C1508 PHI_1 a_32570_158# 0.00164f
C1509 gc[8] DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.33472f
C1510 a_13482_n384# VDD 0.42245f
C1511 Q[7] a_42586_n387# 0
C1512 a_32718_158# PHI_1 0.01804f
C1513 a_5294_158# a_5638_38# 0.57845f
C1514 PHI_1 a_49318_38# 0.01314f
C1515 VDD a_42938_158# 0.01506f
C1516 PHI_1 a_26478_158# 0.01804f
C1517 a_534_n402# PHI_1 0.01733f
C1518 EN DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C1519 Q[9] a_54230_n402# 0.16779f
C1520 gc[5] gc[6] 0.01049f
C1521 a_17774_158# Q[3] 0.01552f
C1522 a_n1094_n387# gc[1] 0
C1523 Q[9] DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C1524 a_13998_158# EN 0.11443f
C1525 a_8102_38# Q[2] 0.25874f
C1526 a_7758_158# DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1527 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN 0.65271f
C1528 a_19722_n384# a_20090_158# 0.00294f
C1529 a_50922_n384# a_51290_158# 0.00294f
C1530 a_51438_158# a_51642_158# 0.01151f
C1531 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_6774_n402# 0.16689f
C1532 a_20442_158# gc[4] 0
C1533 VDD DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C1534 a_57922_n387# a_57678_158# 0.01595f
C1535 a_17258_n384# Q[3] 0.36203f
C1536 EN a_50454_n402# 0.08694f
C1537 gc[8] a_42586_n387# 0
C1538 gc[1] VDD 0.26766f
C1539 a_1370_n387# DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C1540 PHI_2 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C1541 a_24358_38# a_24258_n387# 0
C1542 a_23498_n384# a_23866_n387# 0.00194f
C1543 Q[5] a_25962_n384# 0.00101f
C1544 a_n602_38# PHI_2 0.03207f
C1545 a_17978_158# EN 0.00368f
C1546 a_5294_158# a_4778_n384# 0.30053f
C1547 VDD a_42586_158# 0.00491f
C1548 a_24358_38# a_25494_n402# 0
C1549 PHI_1 a_48458_n384# 0.0533f
C1550 EN a_n1094_158# 0.00101f
C1551 Q[9] a_52903_n425# 0.00241f
C1552 a_16790_n402# Q[3] 0.16779f
C1553 a_n702_n387# gc[1] 0
C1554 gc[7] a_39302_38# 0.01014f
C1555 PHI_1 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.02073f
C1556 a_7242_n384# Q[2] 0.00101f
C1557 a_51438_158# a_51290_158# 0
C1558 a_13998_158# PHI_1 0.01804f
C1559 EN a_44214_n402# 0.08694f
C1560 gc[8] a_46663_n425# 0.00113f
C1561 PHI_2 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C1562 a_18118_38# PHI_2 0.03207f
C1563 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C1564 a_19254_n402# Q[4] 0.00225f
C1565 gc[10] VSS 1.6729f
C1566 Q[10] VSS 1.01569f
C1567 gc[9] VSS 1.65417f
C1568 Q[9] VSS 1.46344f
C1569 gc[8] VSS 1.65417f
C1570 Q[8] VSS 1.46344f
C1571 gc[7] VSS 1.65417f
C1572 Q[7] VSS 1.46344f
C1573 gc[6] VSS 1.65417f
C1574 Q[6] VSS 1.46344f
C1575 gc[5] VSS 1.65417f
C1576 Q[5] VSS 1.46344f
C1577 gc[4] VSS 1.65417f
C1578 Q[4] VSS 1.46344f
C1579 gc[3] VSS 1.65417f
C1580 Q[3] VSS 1.46344f
C1581 gc[2] VSS 1.65417f
C1582 Q[2] VSS 1.46344f
C1583 gc[1] VSS 1.66058f
C1584 EN VSS 28.30377f
C1585 Q[1] VSS 1.46344f
C1586 PHI_2 VSS 19.68128f
C1587 D_in VSS 0.48741f
C1588 PHI_1 VSS 29.6932f
C1589 VDD VSS 0.13498p
C1590 a_59143_n425# VSS 0.0072f
C1591 a_57530_n387# VSS 0.0042f
C1592 a_57922_n387# VSS 0.0095f
C1593 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.77512f
C1594 a_55066_n387# VSS 0.0042f
C1595 a_55458_n387# VSS 0.0095f
C1596 a_58022_38# VSS 0.42076f
C1597 a_57162_n384# VSS 0.53018f
C1598 a_57678_158# VSS 1.13543f
C1599 DFF_2phase_1$1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1600 a_52903_n425# VSS 0.0072f
C1601 a_51290_n387# VSS 0.0042f
C1602 a_51682_n387# VSS 0.0095f
C1603 a_55558_38# VSS 0.42076f
C1604 a_54698_n384# VSS 0.53018f
C1605 a_56694_n402# VSS 1.18728f
C1606 a_55214_158# VSS 1.14251f
C1607 a_54230_n402# VSS 1.18269f
C1608 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1609 a_48826_n387# VSS 0.0042f
C1610 a_49218_n387# VSS 0.0095f
C1611 a_51782_38# VSS 0.42076f
C1612 a_50922_n384# VSS 0.53018f
C1613 a_51438_158# VSS 1.13543f
C1614 DFF_2phase_1$1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1615 a_46663_n425# VSS 0.0072f
C1616 a_45050_n387# VSS 0.0042f
C1617 a_45442_n387# VSS 0.0095f
C1618 a_49318_38# VSS 0.42076f
C1619 a_48458_n384# VSS 0.53018f
C1620 a_50454_n402# VSS 1.18728f
C1621 a_48974_158# VSS 1.14251f
C1622 a_47990_n402# VSS 1.18269f
C1623 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1624 a_42586_n387# VSS 0.0042f
C1625 a_42978_n387# VSS 0.0095f
C1626 a_45542_38# VSS 0.42076f
C1627 a_44682_n384# VSS 0.53018f
C1628 a_45198_158# VSS 1.13543f
C1629 DFF_2phase_1$1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1630 a_40423_n425# VSS 0.0072f
C1631 a_38810_n387# VSS 0.0042f
C1632 a_39202_n387# VSS 0.0095f
C1633 a_43078_38# VSS 0.42076f
C1634 a_42218_n384# VSS 0.53018f
C1635 a_44214_n402# VSS 1.18728f
C1636 a_42734_158# VSS 1.14251f
C1637 a_41750_n402# VSS 1.18269f
C1638 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1639 a_36346_n387# VSS 0.0042f
C1640 a_36738_n387# VSS 0.0095f
C1641 a_39302_38# VSS 0.42076f
C1642 a_38442_n384# VSS 0.53018f
C1643 a_38958_158# VSS 1.13543f
C1644 DFF_2phase_1$1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1645 a_34183_n425# VSS 0.0072f
C1646 a_32570_n387# VSS 0.0042f
C1647 a_32962_n387# VSS 0.0095f
C1648 a_36838_38# VSS 0.42076f
C1649 a_35978_n384# VSS 0.53018f
C1650 a_37974_n402# VSS 1.18728f
C1651 a_36494_158# VSS 1.14251f
C1652 a_35510_n402# VSS 1.18269f
C1653 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1654 a_30106_n387# VSS 0.0042f
C1655 a_30498_n387# VSS 0.0095f
C1656 a_33062_38# VSS 0.42076f
C1657 a_32202_n384# VSS 0.53018f
C1658 a_32718_158# VSS 1.13543f
C1659 DFF_2phase_1$1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1660 a_27943_n425# VSS 0.0072f
C1661 a_26330_n387# VSS 0.0042f
C1662 a_26722_n387# VSS 0.0095f
C1663 a_30598_38# VSS 0.42076f
C1664 a_29738_n384# VSS 0.53018f
C1665 a_31734_n402# VSS 1.18728f
C1666 a_30254_158# VSS 1.14251f
C1667 a_29270_n402# VSS 1.18269f
C1668 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1669 a_23866_n387# VSS 0.0042f
C1670 a_24258_n387# VSS 0.0095f
C1671 a_26822_38# VSS 0.42076f
C1672 a_25962_n384# VSS 0.53018f
C1673 a_26478_158# VSS 1.13543f
C1674 DFF_2phase_1$1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1675 a_21703_n425# VSS 0.0072f
C1676 a_20090_n387# VSS 0.0042f
C1677 a_20482_n387# VSS 0.0095f
C1678 a_24358_38# VSS 0.42076f
C1679 a_23498_n384# VSS 0.53018f
C1680 a_25494_n402# VSS 1.18728f
C1681 a_24014_158# VSS 1.14251f
C1682 a_23030_n402# VSS 1.18269f
C1683 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1684 a_17626_n387# VSS 0.0042f
C1685 a_18018_n387# VSS 0.0095f
C1686 a_20582_38# VSS 0.42076f
C1687 a_19722_n384# VSS 0.53018f
C1688 a_20238_158# VSS 1.13543f
C1689 DFF_2phase_1$1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1690 a_15463_n425# VSS 0.0072f
C1691 a_13850_n387# VSS 0.0042f
C1692 a_14242_n387# VSS 0.0095f
C1693 a_18118_38# VSS 0.42076f
C1694 a_17258_n384# VSS 0.53018f
C1695 a_19254_n402# VSS 1.18728f
C1696 a_17774_158# VSS 1.14251f
C1697 a_16790_n402# VSS 1.18269f
C1698 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1699 a_11386_n387# VSS 0.0042f
C1700 a_11778_n387# VSS 0.0095f
C1701 a_14342_38# VSS 0.42076f
C1702 a_13482_n384# VSS 0.53018f
C1703 a_13998_158# VSS 1.13543f
C1704 DFF_2phase_1$1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1705 a_9223_n425# VSS 0.0072f
C1706 a_7610_n387# VSS 0.0042f
C1707 a_8002_n387# VSS 0.0095f
C1708 a_11878_38# VSS 0.42076f
C1709 a_11018_n384# VSS 0.53018f
C1710 a_13014_n402# VSS 1.18728f
C1711 a_11534_158# VSS 1.14251f
C1712 a_10550_n402# VSS 1.18269f
C1713 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1714 a_5146_n387# VSS 0.0042f
C1715 a_5538_n387# VSS 0.0095f
C1716 a_8102_38# VSS 0.42076f
C1717 a_7242_n384# VSS 0.53018f
C1718 a_7758_158# VSS 1.13543f
C1719 DFF_2phase_1$1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1720 a_2983_n425# VSS 0.0072f
C1721 a_1370_n387# VSS 0.0042f
C1722 a_1762_n387# VSS 0.0095f
C1723 a_5638_38# VSS 0.42076f
C1724 a_4778_n384# VSS 0.53018f
C1725 a_6774_n402# VSS 1.18728f
C1726 a_5294_158# VSS 1.14251f
C1727 a_4310_n402# VSS 1.18269f
C1728 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.76875f
C1729 a_n1094_n387# VSS 0.0042f
C1730 a_n702_n387# VSS 0.0095f
C1731 a_1862_38# VSS 0.42076f
C1732 a_1002_n384# VSS 0.53018f
C1733 a_1518_158# VSS 1.13543f
C1734 DFF_2phase_1$1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C1735 a_n602_38# VSS 0.42076f
C1736 a_n1462_n384# VSS 0.53018f
C1737 a_534_n402# VSS 1.18728f
C1738 a_n946_158# VSS 1.14251f
C1739 a_n1930_n402# VSS 1.19329f
C1740 PHI_2.t4 VSS 0.1095f
C1741 PHI_2.t18 VSS 0.06054f
C1742 PHI_2.n0 VSS 0.10899f
C1743 PHI_2.t15 VSS 0.1095f
C1744 PHI_2.t3 VSS 0.06054f
C1745 PHI_2.n1 VSS 0.10899f
C1746 PHI_2.n2 VSS 1.2589f
C1747 PHI_2.t13 VSS 0.1095f
C1748 PHI_2.t9 VSS 0.06054f
C1749 PHI_2.n3 VSS 0.10899f
C1750 PHI_2.n4 VSS 1.2589f
C1751 PHI_2.t10 VSS 0.1095f
C1752 PHI_2.t1 VSS 0.06054f
C1753 PHI_2.n5 VSS 0.10899f
C1754 PHI_2.n6 VSS 1.2589f
C1755 PHI_2.t16 VSS 0.1095f
C1756 PHI_2.t19 VSS 0.06054f
C1757 PHI_2.n7 VSS 0.10899f
C1758 PHI_2.n8 VSS 1.2589f
C1759 PHI_2.t14 VSS 0.1095f
C1760 PHI_2.t11 VSS 0.06054f
C1761 PHI_2.n9 VSS 0.10899f
C1762 PHI_2.n10 VSS 1.2589f
C1763 PHI_2.t12 VSS 0.1095f
C1764 PHI_2.t17 VSS 0.06054f
C1765 PHI_2.n11 VSS 0.10899f
C1766 PHI_2.n12 VSS 1.2589f
C1767 PHI_2.t5 VSS 0.1095f
C1768 PHI_2.t2 VSS 0.06054f
C1769 PHI_2.n13 VSS 0.10899f
C1770 PHI_2.n14 VSS 1.2589f
C1771 PHI_2.t7 VSS 0.1095f
C1772 PHI_2.t8 VSS 0.06054f
C1773 PHI_2.n15 VSS 0.10899f
C1774 PHI_2.n16 VSS 1.2589f
C1775 PHI_2.t6 VSS 0.1095f
C1776 PHI_2.t0 VSS 0.06054f
C1777 PHI_2.n17 VSS 0.10899f
C1778 PHI_2.n18 VSS 1.2589f
C1779 PHI_1.t7 VSS 0.12714f
C1780 PHI_1.t14 VSS 0.0703f
C1781 PHI_1.n0 VSS 0.1265f
C1782 PHI_1.t4 VSS 0.12714f
C1783 PHI_1.t3 VSS 0.0703f
C1784 PHI_1.n1 VSS 0.1265f
C1785 PHI_1.n2 VSS 1.47113f
C1786 PHI_1.t12 VSS 0.12714f
C1787 PHI_1.t1 VSS 0.0703f
C1788 PHI_1.n3 VSS 0.1265f
C1789 PHI_1.n4 VSS 1.47113f
C1790 PHI_1.t9 VSS 0.12714f
C1791 PHI_1.t15 VSS 0.0703f
C1792 PHI_1.n5 VSS 0.1265f
C1793 PHI_1.n6 VSS 1.47113f
C1794 PHI_1.t6 VSS 0.12714f
C1795 PHI_1.t0 VSS 0.0703f
C1796 PHI_1.n7 VSS 0.1265f
C1797 PHI_1.n8 VSS 1.47113f
C1798 PHI_1.t18 VSS 0.12714f
C1799 PHI_1.t5 VSS 0.0703f
C1800 PHI_1.n9 VSS 0.1265f
C1801 PHI_1.n10 VSS 1.47113f
C1802 PHI_1.t10 VSS 0.12714f
C1803 PHI_1.t11 VSS 0.0703f
C1804 PHI_1.n11 VSS 0.1265f
C1805 PHI_1.n12 VSS 1.47113f
C1806 PHI_1.t2 VSS 0.12714f
C1807 PHI_1.t17 VSS 0.0703f
C1808 PHI_1.n13 VSS 0.1265f
C1809 PHI_1.n14 VSS 1.47113f
C1810 PHI_1.t13 VSS 0.12714f
C1811 PHI_1.t8 VSS 0.0703f
C1812 PHI_1.n15 VSS 0.1265f
C1813 PHI_1.n16 VSS 1.47113f
C1814 PHI_1.t19 VSS 0.12714f
C1815 PHI_1.t16 VSS 0.0703f
C1816 PHI_1.n17 VSS 0.1265f
C1817 PHI_1.n18 VSS 1.47113f
C1818 EN.t17 VSS 0.01373f
C1819 EN.t8 VSS 0.0165f
C1820 EN.n0 VSS 0.01551f
C1821 EN.n1 VSS 0.00498f
C1822 EN.t4 VSS 0.01373f
C1823 EN.t2 VSS 0.0165f
C1824 EN.n2 VSS 0.01551f
C1825 EN.n3 VSS 0.00498f
C1826 EN.t14 VSS 0.01373f
C1827 EN.t9 VSS 0.0165f
C1828 EN.n4 VSS 0.01551f
C1829 EN.n5 VSS 0.00498f
C1830 EN.t18 VSS 0.01373f
C1831 EN.t1 VSS 0.0165f
C1832 EN.n6 VSS 0.01551f
C1833 EN.n7 VSS 0.00498f
C1834 EN.t10 VSS 0.01373f
C1835 EN.t0 VSS 0.0165f
C1836 EN.n8 VSS 0.01551f
C1837 EN.n9 VSS 0.00498f
C1838 EN.t12 VSS 0.01373f
C1839 EN.t13 VSS 0.0165f
C1840 EN.n10 VSS 0.01551f
C1841 EN.n11 VSS 0.00498f
C1842 EN.t15 VSS 0.01373f
C1843 EN.t5 VSS 0.0165f
C1844 EN.n12 VSS 0.01551f
C1845 EN.n13 VSS 0.00498f
C1846 EN.t3 VSS 0.01373f
C1847 EN.t16 VSS 0.0165f
C1848 EN.n14 VSS 0.01551f
C1849 EN.n15 VSS 0.00498f
C1850 EN.t6 VSS 0.01373f
C1851 EN.t11 VSS 0.0165f
C1852 EN.n16 VSS 0.01551f
C1853 EN.n17 VSS 0.00498f
C1854 EN.t19 VSS 0.01373f
C1855 EN.t7 VSS 0.0165f
C1856 EN.n18 VSS 0.01551f
C1857 EN.n19 VSS 0.10138f
C1858 EN.n20 VSS 0.1528f
C1859 EN.n21 VSS 0.1528f
C1860 EN.n22 VSS 0.1528f
C1861 EN.n23 VSS 0.1528f
C1862 EN.n24 VSS 0.1528f
C1863 EN.n25 VSS 0.1528f
C1864 EN.n26 VSS 0.1528f
C1865 EN.n27 VSS 0.1528f
C1866 EN.n28 VSS 0.1528f
C1867 VDD.n0 VSS 0.01993f
C1868 VDD.t215 VSS 0.00346f
C1869 VDD.t114 VSS 0.0017f
C1870 VDD.n1 VSS 0.00736f
C1871 VDD.t286 VSS 0.00432f
C1872 VDD.t178 VSS 0.0023f
C1873 VDD.t230 VSS 0.0023f
C1874 VDD.n2 VSS 0.00491f
C1875 VDD.t180 VSS 0.00873f
C1876 VDD.t265 VSS 0.00752f
C1877 VDD.t238 VSS 0.00742f
C1878 VDD.t106 VSS 0.00858f
C1879 VDD.t113 VSS 0.03957f
C1880 VDD.t214 VSS 0.06454f
C1881 VDD.t285 VSS 0.05303f
C1882 VDD.t213 VSS 0.03617f
C1883 VDD.t126 VSS 0.04563f
C1884 VDD.t229 VSS 0.04563f
C1885 VDD.t177 VSS 0.06495f
C1886 VDD.t179 VSS 0.07101f
C1887 VDD.t264 VSS 0.03186f
C1888 VDD.t237 VSS 0.04666f
C1889 VDD.t105 VSS 0.05005f
C1890 VDD.n3 VSS 0.06545f
C1891 VDD.n4 VSS 0.04726f
C1892 VDD.t206 VSS 0.00346f
C1893 VDD.t251 VSS 0.0017f
C1894 VDD.n5 VSS 0.00736f
C1895 VDD.t143 VSS 0.00432f
C1896 VDD.t339 VSS 0.0023f
C1897 VDD.t8 VSS 0.0023f
C1898 VDD.n6 VSS 0.00491f
C1899 VDD.t337 VSS 0.00873f
C1900 VDD.t250 VSS 0.03957f
C1901 VDD.t205 VSS 0.06454f
C1902 VDD.t142 VSS 0.05303f
C1903 VDD.t204 VSS 0.03617f
C1904 VDD.t267 VSS 0.04563f
C1905 VDD.t7 VSS 0.04563f
C1906 VDD.t338 VSS 0.06495f
C1907 VDD.t336 VSS 0.07502f
C1908 VDD.n7 VSS 0.04706f
C1909 VDD.t57 VSS 0.00346f
C1910 VDD.t110 VSS 0.0017f
C1911 VDD.n8 VSS 0.00736f
C1912 VDD.t78 VSS 0.00432f
C1913 VDD.t133 VSS 0.0023f
C1914 VDD.t26 VSS 0.0023f
C1915 VDD.n9 VSS 0.00491f
C1916 VDD.t131 VSS 0.00873f
C1917 VDD.t119 VSS 0.00752f
C1918 VDD.t188 VSS 0.00742f
C1919 VDD.t316 VSS 0.00858f
C1920 VDD.t109 VSS 0.03957f
C1921 VDD.t56 VSS 0.06454f
C1922 VDD.t77 VSS 0.05303f
C1923 VDD.t55 VSS 0.03617f
C1924 VDD.t318 VSS 0.04563f
C1925 VDD.t25 VSS 0.04563f
C1926 VDD.t132 VSS 0.06495f
C1927 VDD.t130 VSS 0.07101f
C1928 VDD.t118 VSS 0.03186f
C1929 VDD.t187 VSS 0.04666f
C1930 VDD.t315 VSS 0.05005f
C1931 VDD.n10 VSS 0.06545f
C1932 VDD.n11 VSS 0.04726f
C1933 VDD.t314 VSS 0.00346f
C1934 VDD.t184 VSS 0.0017f
C1935 VDD.n12 VSS 0.00736f
C1936 VDD.t276 VSS 0.00432f
C1937 VDD.t168 VSS 0.0023f
C1938 VDD.t279 VSS 0.0023f
C1939 VDD.n13 VSS 0.00491f
C1940 VDD.t166 VSS 0.00873f
C1941 VDD.t183 VSS 0.03957f
C1942 VDD.t313 VSS 0.06454f
C1943 VDD.t275 VSS 0.05303f
C1944 VDD.t312 VSS 0.03617f
C1945 VDD.t272 VSS 0.04563f
C1946 VDD.t278 VSS 0.04563f
C1947 VDD.t167 VSS 0.06495f
C1948 VDD.t165 VSS 0.07502f
C1949 VDD.n14 VSS 0.04706f
C1950 VDD.t72 VSS 0.00346f
C1951 VDD.t259 VSS 0.0017f
C1952 VDD.n15 VSS 0.00736f
C1953 VDD.t48 VSS 0.00432f
C1954 VDD.t60 VSS 0.0023f
C1955 VDD.t108 VSS 0.0023f
C1956 VDD.n16 VSS 0.00491f
C1957 VDD.t62 VSS 0.00873f
C1958 VDD.t248 VSS 0.00752f
C1959 VDD.t232 VSS 0.00742f
C1960 VDD.t284 VSS 0.00858f
C1961 VDD.t258 VSS 0.03957f
C1962 VDD.t71 VSS 0.06454f
C1963 VDD.t47 VSS 0.05303f
C1964 VDD.t70 VSS 0.03617f
C1965 VDD.t317 VSS 0.04563f
C1966 VDD.t107 VSS 0.04563f
C1967 VDD.t59 VSS 0.06495f
C1968 VDD.t61 VSS 0.07101f
C1969 VDD.t247 VSS 0.03186f
C1970 VDD.t231 VSS 0.04666f
C1971 VDD.t283 VSS 0.05005f
C1972 VDD.n17 VSS 0.06545f
C1973 VDD.n18 VSS 0.04726f
C1974 VDD.t289 VSS 0.00346f
C1975 VDD.t253 VSS 0.0017f
C1976 VDD.n19 VSS 0.00736f
C1977 VDD.t141 VSS 0.00432f
C1978 VDD.t85 VSS 0.0023f
C1979 VDD.t89 VSS 0.0023f
C1980 VDD.n20 VSS 0.00491f
C1981 VDD.t83 VSS 0.00873f
C1982 VDD.t252 VSS 0.03957f
C1983 VDD.t288 VSS 0.06454f
C1984 VDD.t140 VSS 0.05303f
C1985 VDD.t290 VSS 0.03617f
C1986 VDD.t38 VSS 0.04563f
C1987 VDD.t88 VSS 0.04563f
C1988 VDD.t84 VSS 0.06495f
C1989 VDD.t82 VSS 0.07502f
C1990 VDD.n21 VSS 0.04706f
C1991 VDD.t154 VSS 0.00346f
C1992 VDD.t326 VSS 0.0017f
C1993 VDD.n22 VSS 0.00736f
C1994 VDD.t164 VSS 0.00432f
C1995 VDD.t137 VSS 0.0023f
C1996 VDD.t139 VSS 0.0023f
C1997 VDD.n23 VSS 0.00491f
C1998 VDD.t135 VSS 0.00873f
C1999 VDD.t91 VSS 0.00752f
C2000 VDD.t257 VSS 0.00742f
C2001 VDD.t192 VSS 0.00858f
C2002 VDD.t325 VSS 0.03957f
C2003 VDD.t153 VSS 0.06454f
C2004 VDD.t163 VSS 0.05303f
C2005 VDD.t152 VSS 0.03617f
C2006 VDD.t49 VSS 0.04563f
C2007 VDD.t138 VSS 0.04563f
C2008 VDD.t136 VSS 0.06495f
C2009 VDD.t134 VSS 0.07101f
C2010 VDD.t90 VSS 0.03186f
C2011 VDD.t256 VSS 0.04666f
C2012 VDD.t191 VSS 0.05005f
C2013 VDD.n24 VSS 0.06545f
C2014 VDD.n25 VSS 0.04726f
C2015 VDD.t282 VSS 0.00346f
C2016 VDD.t145 VSS 0.0017f
C2017 VDD.n26 VSS 0.00736f
C2018 VDD.t324 VSS 0.00432f
C2019 VDD.t160 VSS 0.0023f
C2020 VDD.t40 VSS 0.0023f
C2021 VDD.n27 VSS 0.00491f
C2022 VDD.t162 VSS 0.00873f
C2023 VDD.t144 VSS 0.03957f
C2024 VDD.t281 VSS 0.06454f
C2025 VDD.t323 VSS 0.05303f
C2026 VDD.t280 VSS 0.03617f
C2027 VDD.t117 VSS 0.04563f
C2028 VDD.t39 VSS 0.04563f
C2029 VDD.t159 VSS 0.06495f
C2030 VDD.t161 VSS 0.07502f
C2031 VDD.n28 VSS 0.04706f
C2032 VDD.t42 VSS 0.00346f
C2033 VDD.t330 VSS 0.0017f
C2034 VDD.n29 VSS 0.00736f
C2035 VDD.t170 VSS 0.00432f
C2036 VDD.t271 VSS 0.0023f
C2037 VDD.t81 VSS 0.0023f
C2038 VDD.n30 VSS 0.00491f
C2039 VDD.t269 VSS 0.00873f
C2040 VDD.t322 VSS 0.00752f
C2041 VDD.t186 VSS 0.00742f
C2042 VDD.t307 VSS 0.00858f
C2043 VDD.t329 VSS 0.03957f
C2044 VDD.t41 VSS 0.06454f
C2045 VDD.t169 VSS 0.05303f
C2046 VDD.t43 VSS 0.03617f
C2047 VDD.t266 VSS 0.04563f
C2048 VDD.t80 VSS 0.04563f
C2049 VDD.t270 VSS 0.06495f
C2050 VDD.t268 VSS 0.07101f
C2051 VDD.t321 VSS 0.03186f
C2052 VDD.t185 VSS 0.04666f
C2053 VDD.t306 VSS 0.05005f
C2054 VDD.n31 VSS 0.06545f
C2055 VDD.n32 VSS 0.04726f
C2056 VDD.t76 VSS 0.00346f
C2057 VDD.t182 VSS 0.0017f
C2058 VDD.n33 VSS 0.00736f
C2059 VDD.t320 VSS 0.00432f
C2060 VDD.t37 VSS 0.0023f
C2061 VDD.t102 VSS 0.0023f
C2062 VDD.n34 VSS 0.00491f
C2063 VDD.t35 VSS 0.00873f
C2064 VDD.t181 VSS 0.03957f
C2065 VDD.t75 VSS 0.06454f
C2066 VDD.t319 VSS 0.05303f
C2067 VDD.t74 VSS 0.03617f
C2068 VDD.t73 VSS 0.04563f
C2069 VDD.t101 VSS 0.04563f
C2070 VDD.t36 VSS 0.06495f
C2071 VDD.t34 VSS 0.07502f
C2072 VDD.n35 VSS 0.04706f
C2073 VDD.t53 VSS 0.00346f
C2074 VDD.t217 VSS 0.0017f
C2075 VDD.n36 VSS 0.00736f
C2076 VDD.t295 VSS 0.00432f
C2077 VDD.t98 VSS 0.0023f
C2078 VDD.t172 VSS 0.0023f
C2079 VDD.n37 VSS 0.00491f
C2080 VDD.t96 VSS 0.00873f
C2081 VDD.t194 VSS 0.00752f
C2082 VDD.t244 VSS 0.00742f
C2083 VDD.t87 VSS 0.00858f
C2084 VDD.t216 VSS 0.03957f
C2085 VDD.t52 VSS 0.06454f
C2086 VDD.t294 VSS 0.05303f
C2087 VDD.t54 VSS 0.03617f
C2088 VDD.t333 VSS 0.04563f
C2089 VDD.t171 VSS 0.04563f
C2090 VDD.t97 VSS 0.06495f
C2091 VDD.t95 VSS 0.07101f
C2092 VDD.t193 VSS 0.03186f
C2093 VDD.t243 VSS 0.04666f
C2094 VDD.t86 VSS 0.05005f
C2095 VDD.n38 VSS 0.06545f
C2096 VDD.n39 VSS 0.04726f
C2097 VDD.t129 VSS 0.00346f
C2098 VDD.t240 VSS 0.0017f
C2099 VDD.n40 VSS 0.00736f
C2100 VDD.t196 VSS 0.00432f
C2101 VDD.t305 VSS 0.0023f
C2102 VDD.t21 VSS 0.0023f
C2103 VDD.n41 VSS 0.00491f
C2104 VDD.t303 VSS 0.00873f
C2105 VDD.t239 VSS 0.03957f
C2106 VDD.t128 VSS 0.06454f
C2107 VDD.t195 VSS 0.05303f
C2108 VDD.t127 VSS 0.03617f
C2109 VDD.t249 VSS 0.04563f
C2110 VDD.t20 VSS 0.04563f
C2111 VDD.t304 VSS 0.06495f
C2112 VDD.t302 VSS 0.07502f
C2113 VDD.n42 VSS 0.04706f
C2114 VDD.t23 VSS 0.00346f
C2115 VDD.t261 VSS 0.0017f
C2116 VDD.n43 VSS 0.00736f
C2117 VDD.t274 VSS 0.00432f
C2118 VDD.t123 VSS 0.0023f
C2119 VDD.t208 VSS 0.0023f
C2120 VDD.n44 VSS 0.00491f
C2121 VDD.t125 VSS 0.00873f
C2122 VDD.t299 VSS 0.00752f
C2123 VDD.t236 VSS 0.00742f
C2124 VDD.t311 VSS 0.00858f
C2125 VDD.t260 VSS 0.03957f
C2126 VDD.t22 VSS 0.06454f
C2127 VDD.t273 VSS 0.05303f
C2128 VDD.t24 VSS 0.03617f
C2129 VDD.t287 VSS 0.04563f
C2130 VDD.t207 VSS 0.04563f
C2131 VDD.t122 VSS 0.06495f
C2132 VDD.t124 VSS 0.07101f
C2133 VDD.t298 VSS 0.03186f
C2134 VDD.t235 VSS 0.04666f
C2135 VDD.t310 VSS 0.05005f
C2136 VDD.n45 VSS 0.06545f
C2137 VDD.n46 VSS 0.04726f
C2138 VDD.t11 VSS 0.00346f
C2139 VDD.t228 VSS 0.0017f
C2140 VDD.n47 VSS 0.00736f
C2141 VDD.t297 VSS 0.00432f
C2142 VDD.t222 VSS 0.0023f
C2143 VDD.t100 VSS 0.0023f
C2144 VDD.n48 VSS 0.00491f
C2145 VDD.t224 VSS 0.00873f
C2146 VDD.t227 VSS 0.03957f
C2147 VDD.t10 VSS 0.06454f
C2148 VDD.t296 VSS 0.05303f
C2149 VDD.t9 VSS 0.03617f
C2150 VDD.t293 VSS 0.04563f
C2151 VDD.t99 VSS 0.04563f
C2152 VDD.t221 VSS 0.06495f
C2153 VDD.t223 VSS 0.07502f
C2154 VDD.n49 VSS 0.04706f
C2155 VDD.t46 VSS 0.00346f
C2156 VDD.t328 VSS 0.0017f
C2157 VDD.n50 VSS 0.00736f
C2158 VDD.t64 VSS 0.00432f
C2159 VDD.t174 VSS 0.0023f
C2160 VDD.t212 VSS 0.0023f
C2161 VDD.n51 VSS 0.00491f
C2162 VDD.t176 VSS 0.00873f
C2163 VDD.t2 VSS 0.00752f
C2164 VDD.t263 VSS 0.00742f
C2165 VDD.t121 VSS 0.00858f
C2166 VDD.t327 VSS 0.03957f
C2167 VDD.t45 VSS 0.06454f
C2168 VDD.t63 VSS 0.05303f
C2169 VDD.t44 VSS 0.03617f
C2170 VDD.t277 VSS 0.04563f
C2171 VDD.t211 VSS 0.04563f
C2172 VDD.t173 VSS 0.06495f
C2173 VDD.t175 VSS 0.07101f
C2174 VDD.t1 VSS 0.03186f
C2175 VDD.t262 VSS 0.04666f
C2176 VDD.t120 VSS 0.05005f
C2177 VDD.n52 VSS 0.06545f
C2178 VDD.n53 VSS 0.04726f
C2179 VDD.t202 VSS 0.00346f
C2180 VDD.t147 VSS 0.0017f
C2181 VDD.n54 VSS 0.00736f
C2182 VDD.t4 VSS 0.00432f
C2183 VDD.t151 VSS 0.0023f
C2184 VDD.t332 VSS 0.0023f
C2185 VDD.n55 VSS 0.00491f
C2186 VDD.t149 VSS 0.00873f
C2187 VDD.t146 VSS 0.03957f
C2188 VDD.t201 VSS 0.06454f
C2189 VDD.t3 VSS 0.05303f
C2190 VDD.t203 VSS 0.03617f
C2191 VDD.t0 VSS 0.04563f
C2192 VDD.t331 VSS 0.04563f
C2193 VDD.t150 VSS 0.06495f
C2194 VDD.t148 VSS 0.07502f
C2195 VDD.n56 VSS 0.04706f
C2196 VDD.t220 VSS 0.00346f
C2197 VDD.t116 VSS 0.0017f
C2198 VDD.n57 VSS 0.00736f
C2199 VDD.t69 VSS 0.00432f
C2200 VDD.t200 VSS 0.0023f
C2201 VDD.t6 VSS 0.0023f
C2202 VDD.n58 VSS 0.00491f
C2203 VDD.t198 VSS 0.00873f
C2204 VDD.t292 VSS 0.00752f
C2205 VDD.t234 VSS 0.00742f
C2206 VDD.t51 VSS 0.00858f
C2207 VDD.t115 VSS 0.03957f
C2208 VDD.t219 VSS 0.06454f
C2209 VDD.t68 VSS 0.05303f
C2210 VDD.t218 VSS 0.03617f
C2211 VDD.t158 VSS 0.04563f
C2212 VDD.t5 VSS 0.04563f
C2213 VDD.t199 VSS 0.06495f
C2214 VDD.t197 VSS 0.07101f
C2215 VDD.t291 VSS 0.03186f
C2216 VDD.t233 VSS 0.04666f
C2217 VDD.t50 VSS 0.0507f
C2218 VDD.n59 VSS 0.13062f
C2219 VDD.n60 VSS 0.01984f
C2220 VDD.n61 VSS 0.02095f
C2221 VDD.n62 VSS 0.02849f
C2222 VDD.n63 VSS 0.0448f
C2223 VDD.n64 VSS 0.04042f
C2224 VDD.n65 VSS 0.02783f
C2225 VDD.n66 VSS 0.02501f
C2226 VDD.n67 VSS 0.02939f
C2227 VDD.n68 VSS 0.0448f
C2228 VDD.n69 VSS 0.04042f
C2229 VDD.n70 VSS 0.01969f
C2230 VDD.n71 VSS 0.01993f
C2231 VDD.n72 VSS 0.02496f
C2232 VDD.n73 VSS 0.02302f
C2233 VDD.n74 VSS 0.01984f
C2234 VDD.n75 VSS 0.02095f
C2235 VDD.n76 VSS 0.02849f
C2236 VDD.n77 VSS 0.0448f
C2237 VDD.n78 VSS 0.04042f
C2238 VDD.n79 VSS 0.02783f
C2239 VDD.n80 VSS 0.02501f
C2240 VDD.n81 VSS 0.02939f
C2241 VDD.n82 VSS 0.0448f
C2242 VDD.n83 VSS 0.04042f
C2243 VDD.n84 VSS 0.01969f
C2244 VDD.n85 VSS 0.01993f
C2245 VDD.n86 VSS 0.02496f
C2246 VDD.n87 VSS 0.02302f
C2247 VDD.n88 VSS 0.01984f
C2248 VDD.n89 VSS 0.02095f
C2249 VDD.n90 VSS 0.02849f
C2250 VDD.n91 VSS 0.0448f
C2251 VDD.n92 VSS 0.04042f
C2252 VDD.n93 VSS 0.02783f
C2253 VDD.n94 VSS 0.02501f
C2254 VDD.n95 VSS 0.02939f
C2255 VDD.n96 VSS 0.0448f
C2256 VDD.n97 VSS 0.04042f
C2257 VDD.n98 VSS 0.01969f
C2258 VDD.n99 VSS 0.01993f
C2259 VDD.n100 VSS 0.02496f
C2260 VDD.n101 VSS 0.02302f
C2261 VDD.n102 VSS 0.01984f
C2262 VDD.n103 VSS 0.02095f
C2263 VDD.n104 VSS 0.02849f
C2264 VDD.n105 VSS 0.0448f
C2265 VDD.n106 VSS 0.04042f
C2266 VDD.n107 VSS 0.02783f
C2267 VDD.n108 VSS 0.02501f
C2268 VDD.n109 VSS 0.02939f
C2269 VDD.n110 VSS 0.0448f
C2270 VDD.n111 VSS 0.04042f
C2271 VDD.n112 VSS 0.01969f
C2272 VDD.n113 VSS 0.01993f
C2273 VDD.n114 VSS 0.02496f
C2274 VDD.n115 VSS 0.02302f
C2275 VDD.n116 VSS 0.01984f
C2276 VDD.n117 VSS 0.02095f
C2277 VDD.n118 VSS 0.02849f
C2278 VDD.n119 VSS 0.0448f
C2279 VDD.n120 VSS 0.04042f
C2280 VDD.n121 VSS 0.02783f
C2281 VDD.n122 VSS 0.02501f
C2282 VDD.n123 VSS 0.02939f
C2283 VDD.n124 VSS 0.0448f
C2284 VDD.n125 VSS 0.04042f
C2285 VDD.n126 VSS 0.01969f
C2286 VDD.n127 VSS 0.01993f
C2287 VDD.n128 VSS 0.02496f
C2288 VDD.n129 VSS 0.02302f
C2289 VDD.n130 VSS 0.01984f
C2290 VDD.n131 VSS 0.02095f
C2291 VDD.n132 VSS 0.02849f
C2292 VDD.n133 VSS 0.0448f
C2293 VDD.n134 VSS 0.04042f
C2294 VDD.n135 VSS 0.02783f
C2295 VDD.n136 VSS 0.02501f
C2296 VDD.n137 VSS 0.02939f
C2297 VDD.n138 VSS 0.0448f
C2298 VDD.n139 VSS 0.04042f
C2299 VDD.n140 VSS 0.01969f
C2300 VDD.n141 VSS 0.01993f
C2301 VDD.n142 VSS 0.02496f
C2302 VDD.n143 VSS 0.02302f
C2303 VDD.n144 VSS 0.01984f
C2304 VDD.n145 VSS 0.02095f
C2305 VDD.n146 VSS 0.02849f
C2306 VDD.n147 VSS 0.0448f
C2307 VDD.n148 VSS 0.04042f
C2308 VDD.n149 VSS 0.02783f
C2309 VDD.n150 VSS 0.02501f
C2310 VDD.n151 VSS 0.02939f
C2311 VDD.n152 VSS 0.0448f
C2312 VDD.n153 VSS 0.04042f
C2313 VDD.n154 VSS 0.01969f
C2314 VDD.n155 VSS 0.01993f
C2315 VDD.n156 VSS 0.02496f
C2316 VDD.n157 VSS 0.02302f
C2317 VDD.n158 VSS 0.01984f
C2318 VDD.n159 VSS 0.02095f
C2319 VDD.n160 VSS 0.02849f
C2320 VDD.n161 VSS 0.0448f
C2321 VDD.n162 VSS 0.04042f
C2322 VDD.n163 VSS 0.02783f
C2323 VDD.n164 VSS 0.02501f
C2324 VDD.n165 VSS 0.02939f
C2325 VDD.n166 VSS 0.0448f
C2326 VDD.n167 VSS 0.04042f
C2327 VDD.n168 VSS 0.01969f
C2328 VDD.n169 VSS 0.01993f
C2329 VDD.n170 VSS 0.02496f
C2330 VDD.n171 VSS 0.02302f
C2331 VDD.n172 VSS 0.01984f
C2332 VDD.n173 VSS 0.02095f
C2333 VDD.n174 VSS 0.02849f
C2334 VDD.n175 VSS 0.0448f
C2335 VDD.n176 VSS 0.04042f
C2336 VDD.n177 VSS 0.02783f
C2337 VDD.t17 VSS 0.00873f
C2338 VDD.t19 VSS 0.0023f
C2339 VDD.t309 VSS 0.0023f
C2340 VDD.n178 VSS 0.00491f
C2341 VDD.t190 VSS 0.00432f
C2342 VDD.t157 VSS 0.00346f
C2343 VDD.t242 VSS 0.0017f
C2344 VDD.n179 VSS 0.00736f
C2345 VDD.n180 VSS 0.01969f
C2346 VDD.n181 VSS 0.04042f
C2347 VDD.n182 VSS 0.0448f
C2348 VDD.n183 VSS 0.02939f
C2349 VDD.n184 VSS 0.02501f
C2350 VDD.n185 VSS 0.04706f
C2351 VDD.t16 VSS 0.07502f
C2352 VDD.t18 VSS 0.06495f
C2353 VDD.t308 VSS 0.04563f
C2354 VDD.t79 VSS 0.04563f
C2355 VDD.t155 VSS 0.03617f
C2356 VDD.t189 VSS 0.05303f
C2357 VDD.t156 VSS 0.06454f
C2358 VDD.t241 VSS 0.03957f
C2359 VDD.n186 VSS 0.04726f
C2360 VDD.n187 VSS 0.06545f
C2361 VDD.t104 VSS 0.00858f
C2362 VDD.t246 VSS 0.00742f
C2363 VDD.t226 VSS 0.00752f
C2364 VDD.t13 VSS 0.00873f
C2365 VDD.t15 VSS 0.0023f
C2366 VDD.t335 VSS 0.0023f
C2367 VDD.n188 VSS 0.00491f
C2368 VDD.t301 VSS 0.00432f
C2369 VDD.t67 VSS 0.00346f
C2370 VDD.t112 VSS 0.0017f
C2371 VDD.n189 VSS 0.00736f
C2372 VDD.t103 VSS 0.05005f
C2373 VDD.t245 VSS 0.04666f
C2374 VDD.t225 VSS 0.03186f
C2375 VDD.t12 VSS 0.07101f
C2376 VDD.t14 VSS 0.06495f
C2377 VDD.t334 VSS 0.04563f
C2378 VDD.t94 VSS 0.04563f
C2379 VDD.t65 VSS 0.03617f
C2380 VDD.t300 VSS 0.05303f
C2381 VDD.t66 VSS 0.06454f
C2382 VDD.t111 VSS 0.03957f
C2383 VDD.n190 VSS 0.04706f
C2384 VDD.t33 VSS 0.00873f
C2385 VDD.t31 VSS 0.0023f
C2386 VDD.t93 VSS 0.0023f
C2387 VDD.n191 VSS 0.00491f
C2388 VDD.t210 VSS 0.00432f
C2389 VDD.t28 VSS 0.00346f
C2390 VDD.t255 VSS 0.0017f
C2391 VDD.n192 VSS 0.00736f
C2392 VDD.t32 VSS 0.07502f
C2393 VDD.t30 VSS 0.06495f
C2394 VDD.t92 VSS 0.04563f
C2395 VDD.t58 VSS 0.04563f
C2396 VDD.t29 VSS 0.03617f
C2397 VDD.t209 VSS 0.05303f
C2398 VDD.t27 VSS 0.06454f
C2399 VDD.t254 VSS 0.03957f
C2400 VDD.n193 VSS 0.07496f
C2401 VDD.n194 VSS 0.01969f
C2402 VDD.n195 VSS 0.04042f
C2403 VDD.n196 VSS 0.0448f
C2404 VDD.n197 VSS 0.02939f
C2405 VDD.n198 VSS 0.02501f
C2406 VDD.n199 VSS 0.02783f
C2407 VDD.n200 VSS 0.04042f
C2408 VDD.n201 VSS 0.0448f
C2409 VDD.n202 VSS 0.02849f
C2410 VDD.n203 VSS 0.02095f
C2411 VDD.n204 VSS 0.01984f
C2412 VDD.n205 VSS 0.02302f
C2413 VDD.n206 VSS 0.02496f
.ends

