magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l36d0 >>
<< l38d0 >>
<< l42d0 >>
<< end >>
