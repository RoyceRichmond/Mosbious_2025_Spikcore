* Extracted by KLayout with GF180 LVS runset on : 12/08/2025 02:36

.SUBCKT DFF_2phase_1 VSS E|PHI_2 D|Q|out_m Q VDD D E|PHI_1 gf180mcu_gnd
M$1 VDD \$26 D|Q|out_m VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$2 \$37 D VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$3 \$26 \$23 \$37 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U PD=1.52U
M$4 \$26 \$24 \$39 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$5 VDD \$27 \$39 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$6 \$27 \$26 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$7 VDD E|PHI_2 \$2 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$8 \$4 \$2 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U PD=2.88U
M$9 VDD E|PHI_1 \$23 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$10 \$24 \$23 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$11 \$20 D|Q|out_m VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$12 \$6 \$2 \$20 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U PD=1.52U
M$13 \$6 \$4 \$21 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U PD=1.52U
M$14 VDD \$7 \$21 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$15 \$7 \$6 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$16 VDD \$6 Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$17 VSS \$26 D|Q|out_m gf180mcu_gnd nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$18 \$29 D VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$19 \$26 \$24 \$29 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$20 \$35 \$23 \$26 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$21 VSS \$27 \$35 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$22 \$27 \$26 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$23 VSS E|PHI_1 \$23 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.3476P
+ AD=0.263P PS=2.46U PD=1.49U
M$24 \$24 \$23 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$25 \$11 D|Q|out_m VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.308P
+ AD=0.084P PS=2.28U PD=0.94U
M$26 \$6 \$4 \$11 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$27 \$13 \$2 \$6 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$28 VSS \$7 \$13 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$29 \$7 \$6 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$30 VSS E|PHI_2 \$2 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$31 \$4 \$2 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$32 VSS \$6 Q gf180mcu_gnd nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
.ENDS DFF_2phase_1
