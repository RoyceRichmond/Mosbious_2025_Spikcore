magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l33d0 >>
<< l34d0 >>
<< l30d0 >>
<< l22d0 >>
<< l31d0 >>
<< l49d0 >>
<< l110d5 >>
<< labels >>
rlabel l34d10 -0.033 0.215 -0.033 0.215 0 
rlabel l34d10 0.133 0.215 0.133 0.215 0 
rlabel l34d10 -0.17 0.215 -0.17 0.215 0 
<< end >>
