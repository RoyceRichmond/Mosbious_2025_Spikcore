** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/pex/AH_neuron/AH_neuron_pex.sch
**.subckt AH_neuron_pex
V1 net2 vss 3.3
I0 vdd net1 PULSE(0 1000p 1u 10n 10n 1u 5u)
R1 vdd net2 10 m=1
R2 vout vss 250k m=1
Vdd_c1 net1 vmem 0
.save i(vdd_c1)
V2 net3 GND 0.49
R3 v_bias net3 10 m=1
V3 vss GND 0
x1 vdd vmem vout vss v_bias AH_neuron
**** begin user architecture code


.option method=gear seed=12
.include /foss/designs/Mosbious_2025_Spikcore/designs/pex/AH_neuron/AH_neuron_pex.spice
.tran 100n 5m
.param vd_v=3.3
.save allcurrents
.options save currents
.control
	reset
	save all
        run
        write AH_neuron_pex.raw
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
