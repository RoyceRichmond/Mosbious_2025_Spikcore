* NGSPICE file created from TG_bootstrapped.ext - technology: gf180mcuD
.subckt TG_bootstrapped_pex vdd vss clk nclk vin vout
X0 vout.t21 a_5673_n171# a_5757_n39.t5 vss.t24 nfet_03v3 ad=2.38815p pd=9.05u as=1.0179p ps=4.435u w=3.915u l=0.42u
X1 a_5757_n39.t4 a_5673_n171# vout.t20 vss.t23 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X2 a_5381_1389.t19 a_5297_1329.t4 vout.t24 vdd.t22 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X3 a_8039_2775# a_5944_2887# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X4 vin.t3 clk.t0 a_8039_2775# vss.t25 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X5 a_5381_1389.t18 a_5297_1329.t5 vout.t32 vdd.t21 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X6 vout.t2 a_5297_1329.t6 a_5381_1389.t17 vdd.t20 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X7 vout.t5 a_5297_1329.t7 a_5381_1389.t16 vdd.t19 pfet_03v3 ad=2.028p pd=7.54u as=0.8112p ps=3.64u w=3.12u l=0.42u
X8 a_5381_1389.t15 a_5297_1329.t8 vout.t22 vdd.t18 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X9 a_5381_1389.t14 a_5297_1329.t9 vout.t3 vdd.t17 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X10 vss.t2 nclk.t0 a_5673_n171# vss.t1 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X11 vout.t35 a_5297_1329.t10 a_5381_1389.t13 vdd.t16 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X12 a_5381_1389.t12 a_5297_1329.t11 vout.t0 vdd.t15 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X13 a_5381_1389.t11 a_5297_1329.t12 vout.t1 vdd.t14 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X14 a_8034_n1134# nclk.t1 vss.t5 vss.t4 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X15 vin.t1 nclk.t2 a_8034_n1134# vdd.t23 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X16 a_5757_n39.t2 a_5673_n171# vout.t19 vss.t22 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X17 vout.t18 a_5673_n171# a_5757_n39.t15 vss.t21 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X18 vout.t17 a_5673_n171# a_5757_n39.t14 vss.t20 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X19 vout.t16 a_5673_n171# a_5757_n39.t13 vss.t19 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X20 vdd.t27 clk.t1 a_5297_1329.t2 vdd.t26 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X21 a_5757_n39.t12 a_5673_n171# vout.t15 vss.t18 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X22 a_5904_n1280# clk.t2 vss.t8 vss.t7 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X23 a_5297_1329.t1 nclk.t3 a_5944_2887# vdd.t1 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X24 a_5673_n171# nclk.t4 a_5904_n1280# vdd.t0 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X25 a_5381_1389.t10 a_5297_1329.t13 vout.t30 vdd.t13 pfet_03v3 ad=0.8112p pd=3.64u as=2.028p ps=7.54u w=3.12u l=0.42u
X26 vout.t26 a_5297_1329.t14 a_5381_1389.t9 vdd.t12 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X27 vout.t27 a_5297_1329.t15 a_5381_1389.t8 vdd.t11 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X28 vout.t25 a_5297_1329.t16 a_5381_1389.t7 vdd.t10 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X29 a_5381_1389.t6 a_5297_1329.t17 vout.t33 vdd.t9 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X30 a_8034_n1134# a_5904_n1280# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X31 vin.t0 nclk.t5 a_8039_2775# vdd.t2 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X32 vdd.t28 nclk.t6 a_5297_1329.t3 vss.t26 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X33 a_5297_1329.t0 clk.t3 a_5944_2887# vss.t0 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X34 a_5757_n39.t11 a_5673_n171# vout.t14 vss.t17 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X35 vss.t27 clk.t4 a_5673_n171# vdd.t31 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X36 a_5757_n39.t10 a_5673_n171# vout.t13 vss.t16 nfet_03v3 ad=1.0179p pd=4.435u as=2.38815p ps=9.05u w=3.915u l=0.42u
X37 a_5757_n39.t1 a_5673_n171# vout.t12 vss.t15 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X38 vout.t11 a_5673_n171# a_5757_n39.t0 vss.t14 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X39 vdd.t30 nclk.t7 a_8039_2775# vdd.t29 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X40 vout.t10 a_5673_n171# a_5757_n39.t9 vss.t13 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X41 vout.t29 a_5297_1329.t18 a_5381_1389.t5 vdd.t8 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X42 a_5381_1389.t4 a_5297_1329.t19 vout.t28 vdd.t7 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X43 a_5944_2887# clk.t5 vdd.t25 vdd.t24 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X44 vout.t31 a_5297_1329.t20 a_5381_1389.t3 vdd.t6 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X45 vout.t23 a_5297_1329.t21 a_5381_1389.t2 vdd.t5 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X46 vout.t4 a_5297_1329.t22 a_5381_1389.t1 vdd.t4 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X47 a_5381_1389.t0 a_5297_1329.t23 vout.t34 vdd.t3 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X48 vout.t9 a_5673_n171# a_5757_n39.t8 vss.t12 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X49 vin.t2 clk.t6 a_8034_n1134# vss.t3 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X50 vout.t8 a_5673_n171# a_5757_n39.t7 vss.t11 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X51 a_5757_n39.t6 a_5673_n171# vout.t7 vss.t10 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X52 a_5757_n39.t3 a_5673_n171# vout.t6 vss.t9 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X53 a_5673_n171# clk.t7 a_5904_n1280# vss.t6 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
R0 a_5757_n39.n12 a_5757_n39.n0 1.91808
R1 a_5757_n39.n3 a_5757_n39.n1 1.91808
R2 a_5757_n39.n11 a_5757_n39.n10 1.86521
R3 a_5757_n39.n9 a_5757_n39.n8 1.86521
R4 a_5757_n39.n7 a_5757_n39.n6 1.86521
R5 a_5757_n39.n5 a_5757_n39.n4 1.86521
R6 a_5757_n39.n3 a_5757_n39.n2 1.86521
R7 a_5757_n39.n13 a_5757_n39.n12 1.86452
R8 a_5757_n39.n1 a_5757_n39.t7 0.418891
R9 a_5757_n39.n1 a_5757_n39.t10 0.418891
R10 a_5757_n39.n2 a_5757_n39.t14 0.418891
R11 a_5757_n39.n2 a_5757_n39.t4 0.418891
R12 a_5757_n39.n4 a_5757_n39.t8 0.418891
R13 a_5757_n39.n4 a_5757_n39.t1 0.418891
R14 a_5757_n39.n6 a_5757_n39.t13 0.418891
R15 a_5757_n39.n6 a_5757_n39.t2 0.418891
R16 a_5757_n39.n8 a_5757_n39.t9 0.418891
R17 a_5757_n39.n8 a_5757_n39.t12 0.418891
R18 a_5757_n39.n10 a_5757_n39.t15 0.418891
R19 a_5757_n39.n10 a_5757_n39.t6 0.418891
R20 a_5757_n39.n0 a_5757_n39.t5 0.418891
R21 a_5757_n39.n0 a_5757_n39.t3 0.418891
R22 a_5757_n39.t0 a_5757_n39.n13 0.418891
R23 a_5757_n39.n13 a_5757_n39.t11 0.418891
R24 a_5757_n39.n12 a_5757_n39.n11 0.053375
R25 a_5757_n39.n11 a_5757_n39.n9 0.053375
R26 a_5757_n39.n9 a_5757_n39.n7 0.053375
R27 a_5757_n39.n7 a_5757_n39.n5 0.053375
R28 a_5757_n39.n5 a_5757_n39.n3 0.053375
R29 vout.n1 vout.t5 2.56303
R30 vout.n28 vout.t30 2.56303
R31 vout.n29 vout.n26 2.31025
R32 vout.n31 vout.n26 2.2505
R33 vout.n33 vout.n32 2.2505
R34 vout.n35 vout.n34 2.2505
R35 vout.n36 vout.n20 2.2505
R36 vout.n39 vout.n38 2.2505
R37 vout.n40 vout.n19 2.2505
R38 vout.n42 vout.n41 2.2505
R39 vout.n44 vout.n16 2.2505
R40 vout.n46 vout.n45 2.2505
R41 vout.n48 vout.n47 2.2505
R42 vout.n49 vout.n10 2.2505
R43 vout.n52 vout.n51 2.2505
R44 vout.n53 vout.n9 2.2505
R45 vout.n55 vout.n54 2.2505
R46 vout.n57 vout.n6 2.2505
R47 vout.n59 vout.n58 2.2505
R48 vout.n61 vout.n60 2.2505
R49 vout.n62 vout.n0 2.2505
R50 vout.n65 vout.n64 2.2505
R51 vout.n28 vout.t13 2.24523
R52 vout.n1 vout.t21 2.24523
R53 vout.n5 vout.n4 1.60155
R54 vout.n56 vout.n8 1.60155
R55 vout.n50 vout.n12 1.60155
R56 vout.n15 vout.n14 1.60155
R57 vout.n43 vout.n18 1.60155
R58 vout.n37 vout.n22 1.60155
R59 vout.n25 vout.n24 1.60155
R60 vout.n63 vout.n2 1.47822
R61 vout.n5 vout.n3 1.47822
R62 vout.n56 vout.n7 1.47822
R63 vout.n50 vout.n11 1.47822
R64 vout.n15 vout.n13 1.47822
R65 vout.n43 vout.n17 1.47822
R66 vout.n37 vout.n21 1.47822
R67 vout.n25 vout.n23 1.47822
R68 vout.n30 vout.n27 1.47822
R69 vout vout.n65 1.02411
R70 vout.n2 vout.t24 0.583833
R71 vout.n2 vout.t29 0.583833
R72 vout.n3 vout.t1 0.583833
R73 vout.n3 vout.t4 0.583833
R74 vout.n7 vout.t0 0.583833
R75 vout.n7 vout.t2 0.583833
R76 vout.n11 vout.t28 0.583833
R77 vout.n11 vout.t25 0.583833
R78 vout.n13 vout.t3 0.583833
R79 vout.n13 vout.t27 0.583833
R80 vout.n17 vout.t22 0.583833
R81 vout.n17 vout.t23 0.583833
R82 vout.n21 vout.t33 0.583833
R83 vout.n21 vout.t35 0.583833
R84 vout.n23 vout.t34 0.583833
R85 vout.n23 vout.t26 0.583833
R86 vout.n27 vout.t32 0.583833
R87 vout.n27 vout.t31 0.583833
R88 vout.n4 vout.t6 0.418891
R89 vout.n4 vout.t11 0.418891
R90 vout.n8 vout.t14 0.418891
R91 vout.n8 vout.t18 0.418891
R92 vout.n12 vout.t7 0.418891
R93 vout.n12 vout.t10 0.418891
R94 vout.n14 vout.t15 0.418891
R95 vout.n14 vout.t16 0.418891
R96 vout.n18 vout.t19 0.418891
R97 vout.n18 vout.t9 0.418891
R98 vout.n22 vout.t12 0.418891
R99 vout.n22 vout.t17 0.418891
R100 vout.n24 vout.t20 0.418891
R101 vout.n24 vout.t8 0.418891
R102 vout.n62 vout.n61 0.0605
R103 vout.n58 vout.n57 0.0605
R104 vout.n55 vout.n9 0.0605
R105 vout.n51 vout.n9 0.0605
R106 vout.n49 vout.n48 0.0605
R107 vout.n45 vout.n44 0.0605
R108 vout.n42 vout.n19 0.0605
R109 vout.n38 vout.n19 0.0605
R110 vout.n36 vout.n35 0.0605
R111 vout.n32 vout.n31 0.0605
R112 vout.n65 vout.n0 0.060251
R113 vout.n60 vout.n0 0.060251
R114 vout.n60 vout.n59 0.060251
R115 vout.n59 vout.n6 0.060251
R116 vout.n54 vout.n6 0.060251
R117 vout.n54 vout.n53 0.060251
R118 vout.n53 vout.n52 0.060251
R119 vout.n52 vout.n10 0.060251
R120 vout.n47 vout.n10 0.060251
R121 vout.n47 vout.n46 0.060251
R122 vout.n46 vout.n16 0.060251
R123 vout.n41 vout.n16 0.060251
R124 vout.n41 vout.n40 0.060251
R125 vout.n40 vout.n39 0.060251
R126 vout.n39 vout.n20 0.060251
R127 vout.n34 vout.n20 0.060251
R128 vout.n34 vout.n33 0.060251
R129 vout.n33 vout.n26 0.060251
R130 vout.n63 vout.n62 0.05525
R131 vout.n31 vout.n30 0.05375
R132 vout.n50 vout.n49 0.05225
R133 vout.n44 vout.n43 0.05075
R134 vout.n37 vout.n36 0.04925
R135 vout.n57 vout.n56 0.04775
R136 vout.n58 vout.n5 0.03425
R137 vout.n35 vout.n25 0.03275
R138 vout.n45 vout.n15 0.03125
R139 vout.n48 vout.n15 0.02975
R140 vout.n32 vout.n25 0.02825
R141 vout.n61 vout.n5 0.02675
R142 vout.n56 vout.n55 0.01325
R143 vout.n38 vout.n37 0.01175
R144 vout.n43 vout.n42 0.01025
R145 vout.n51 vout.n50 0.00875
R146 vout.n30 vout.n29 0.00725
R147 vout.n64 vout.n1 0.00575
R148 vout.n64 vout.n63 0.00575
R149 vout.n29 vout.n28 0.00425
R150 vss.n14 vss.n13 28130.3
R151 vss.n13 vss.n3 3658.85
R152 vss.n15 vss.n14 3473.68
R153 vss.n14 vss.t0 2794.63
R154 vss.n13 vss.t4 2578.99
R155 vss.t3 vss.t1 1060.25
R156 vss.t25 vss.t26 920.038
R157 vss.n12 vss.t6 541.668
R158 vss.t1 vss.n20 480.928
R159 vss.n20 vss.t6 480.928
R160 vss.n23 vss.t3 470.882
R161 vss.t26 vss.n2 416.243
R162 vss.t0 vss.n2 416.243
R163 vss.n3 vss.t25 406.25
R164 vss.n24 vss.t24 358.844
R165 vss.t9 vss.t24 319.728
R166 vss.t14 vss.t9 319.728
R167 vss.t17 vss.t14 319.728
R168 vss.t21 vss.t17 319.728
R169 vss.t10 vss.t21 319.728
R170 vss.t13 vss.t10 319.728
R171 vss.t18 vss.t13 319.728
R172 vss.t19 vss.t18 319.728
R173 vss.t22 vss.t19 319.728
R174 vss.t12 vss.t22 319.728
R175 vss.t15 vss.t12 319.728
R176 vss.t20 vss.t15 319.728
R177 vss.n24 vss.n23 301.611
R178 vss.t4 vss.n7 175.298
R179 vss.t11 vss.t23 131.823
R180 vss.n12 vss.t20 122.45
R181 vss.t16 vss.t7 112.891
R182 vss.n25 vss.n7 86.9476
R183 vss.t23 vss.n12 81.3381
R184 vss.n15 vss.t16 62.4061
R185 vss.n25 vss.n24 37.1634
R186 vss.n28 vss.n3 19.8888
R187 vss.n23 vss.n22 19.6851
R188 vss.t7 vss.t11 18.9325
R189 vss.n17 vss.n16 11.0839
R190 vss.n16 vss.t8 10.8815
R191 vss.n21 vss.t5 10.877
R192 vss.n21 vss.n7 10.4837
R193 vss.n16 vss.n15 10.4793
R194 vss.n5 vss.t2 9.6559
R195 vss.n22 vss.n21 9.22213
R196 vss.n33 vss.n32 4.59325
R197 vss.n10 vss.n8 4.59325
R198 vss.n31 vss.n30 4.5005
R199 vss.n19 vss.n18 4.5005
R200 vss.n11 vss.n9 4.5005
R201 vss.n18 vss.n17 4.5005
R202 vss.n1 vss.n0 4.5005
R203 vss.n30 vss.n29 4.5005
R204 vss.n26 vss.n25 3.80854
R205 vss.n5 vss.t27 3.71674
R206 vss.n6 vss.n5 2.94978
R207 vss.n32 vss.n31 2.20487
R208 vss.n19 vss.n8 2.20487
R209 vss.n26 vss.n6 1.34213
R210 vss.n27 vss.n4 1.02307
R211 vss.n28 vss.n27 0.918196
R212 vss vss.n33 0.60333
R213 vss.n22 vss.n4 0.4415
R214 vss.n31 vss.n2 0.298561
R215 vss.n29 vss.n28 0.280052
R216 vss.n20 vss.n19 0.271533
R217 vss.n27 vss.n26 0.201851
R218 vss.n30 vss.n1 0.188872
R219 vss.n18 vss.n9 0.188872
R220 vss.n22 vss.n6 0.176
R221 vss.n10 vss.n4 0.0973229
R222 vss.n32 vss.n1 0.0932551
R223 vss.n9 vss.n8 0.0932551
R224 vss.n29 vss.n0 0.0387075
R225 vss.n33 vss.n0 0.0387075
R226 vss.n11 vss.n10 0.0116647
R227 vss.n17 vss.n11 0.0116647
R228 a_5297_1329.n3 a_5297_1329.t13 43.8541
R229 a_5297_1329.n14 a_5297_1329.t7 43.8541
R230 a_5297_1329.n3 a_5297_1329.t20 43.6315
R231 a_5297_1329.n4 a_5297_1329.t5 43.6315
R232 a_5297_1329.n5 a_5297_1329.t14 43.6315
R233 a_5297_1329.n6 a_5297_1329.t23 43.6315
R234 a_5297_1329.n7 a_5297_1329.t10 43.6315
R235 a_5297_1329.n8 a_5297_1329.t17 43.6315
R236 a_5297_1329.n9 a_5297_1329.t21 43.6315
R237 a_5297_1329.n12 a_5297_1329.t8 43.6315
R238 a_5297_1329.n11 a_5297_1329.t15 43.6315
R239 a_5297_1329.n22 a_5297_1329.t9 43.6315
R240 a_5297_1329.n21 a_5297_1329.t16 43.6315
R241 a_5297_1329.n20 a_5297_1329.t19 43.6315
R242 a_5297_1329.n19 a_5297_1329.t6 43.6315
R243 a_5297_1329.n18 a_5297_1329.t11 43.6315
R244 a_5297_1329.n17 a_5297_1329.t22 43.6315
R245 a_5297_1329.n16 a_5297_1329.t12 43.6315
R246 a_5297_1329.n15 a_5297_1329.t18 43.6315
R247 a_5297_1329.n14 a_5297_1329.t4 43.6315
R248 a_5297_1329.n26 a_5297_1329.t3 9.65161
R249 a_5297_1329.t0 a_5297_1329.n32 9.65118
R250 a_5297_1329.n24 a_5297_1329.n10 9.0005
R251 a_5297_1329.n24 a_5297_1329.n13 9.0005
R252 a_5297_1329.n24 a_5297_1329.n2 9.0005
R253 a_5297_1329.n24 a_5297_1329.n23 9.0005
R254 a_5297_1329.n29 a_5297_1329.n27 4.5005
R255 a_5297_1329.n30 a_5297_1329.n25 4.5005
R256 a_5297_1329.n31 a_5297_1329.n30 4.5005
R257 a_5297_1329.n30 a_5297_1329.n29 4.5005
R258 a_5297_1329.n32 a_5297_1329.t1 3.70851
R259 a_5297_1329.n26 a_5297_1329.t2 3.7081
R260 a_5297_1329.n28 a_5297_1329.n1 2.24497
R261 a_5297_1329.n27 a_5297_1329.n0 2.24204
R262 a_5297_1329.n29 a_5297_1329.n26 1.04096
R263 a_5297_1329.n32 a_5297_1329.n31 1.03826
R264 a_5297_1329.n9 a_5297_1329.n8 0.223132
R265 a_5297_1329.n8 a_5297_1329.n7 0.223132
R266 a_5297_1329.n7 a_5297_1329.n6 0.223132
R267 a_5297_1329.n6 a_5297_1329.n5 0.223132
R268 a_5297_1329.n5 a_5297_1329.n4 0.223132
R269 a_5297_1329.n4 a_5297_1329.n3 0.223132
R270 a_5297_1329.n15 a_5297_1329.n14 0.223132
R271 a_5297_1329.n16 a_5297_1329.n15 0.223132
R272 a_5297_1329.n17 a_5297_1329.n16 0.223132
R273 a_5297_1329.n18 a_5297_1329.n17 0.223132
R274 a_5297_1329.n19 a_5297_1329.n18 0.223132
R275 a_5297_1329.n20 a_5297_1329.n19 0.223132
R276 a_5297_1329.n21 a_5297_1329.n20 0.223132
R277 a_5297_1329.n23 a_5297_1329.n22 0.153263
R278 a_5297_1329.n11 a_5297_1329.n2 0.139053
R279 a_5297_1329.n13 a_5297_1329.n12 0.124842
R280 a_5297_1329.n30 a_5297_1329.n24 0.114452
R281 a_5297_1329.n10 a_5297_1329.n9 0.110632
R282 a_5297_1329.n12 a_5297_1329.n10 0.108263
R283 a_5297_1329.n13 a_5297_1329.n11 0.0940526
R284 a_5297_1329.n22 a_5297_1329.n2 0.0798421
R285 a_5297_1329.n23 a_5297_1329.n21 0.0656316
R286 a_5297_1329.n29 a_5297_1329.n28 0.0365
R287 a_5297_1329.n28 a_5297_1329.n25 0.0365
R288 a_5297_1329.n31 a_5297_1329.n0 0.0189283
R289 a_5297_1329.n25 a_5297_1329.n0 0.0189283
R290 a_5297_1329.n30 a_5297_1329.n1 0.0130643
R291 a_5297_1329.n27 a_5297_1329.n1 0.0130643
R292 a_5381_1389.n2 a_5381_1389.n0 2.12064
R293 a_5381_1389.n16 a_5381_1389.n15 2.12064
R294 a_5381_1389.n2 a_5381_1389.n1 2.05296
R295 a_5381_1389.n4 a_5381_1389.n3 2.05296
R296 a_5381_1389.n6 a_5381_1389.n5 2.05296
R297 a_5381_1389.n8 a_5381_1389.n7 2.05296
R298 a_5381_1389.n10 a_5381_1389.n9 2.05296
R299 a_5381_1389.n12 a_5381_1389.n11 2.05296
R300 a_5381_1389.n14 a_5381_1389.n13 2.05296
R301 a_5381_1389.n17 a_5381_1389.n16 2.05239
R302 a_5381_1389.n15 a_5381_1389.t3 0.583833
R303 a_5381_1389.n15 a_5381_1389.t10 0.583833
R304 a_5381_1389.n13 a_5381_1389.t13 0.583833
R305 a_5381_1389.n13 a_5381_1389.t0 0.583833
R306 a_5381_1389.n11 a_5381_1389.t2 0.583833
R307 a_5381_1389.n11 a_5381_1389.t6 0.583833
R308 a_5381_1389.n9 a_5381_1389.t8 0.583833
R309 a_5381_1389.n9 a_5381_1389.t15 0.583833
R310 a_5381_1389.n7 a_5381_1389.t7 0.583833
R311 a_5381_1389.n7 a_5381_1389.t14 0.583833
R312 a_5381_1389.n5 a_5381_1389.t17 0.583833
R313 a_5381_1389.n5 a_5381_1389.t4 0.583833
R314 a_5381_1389.n3 a_5381_1389.t1 0.583833
R315 a_5381_1389.n3 a_5381_1389.t12 0.583833
R316 a_5381_1389.n1 a_5381_1389.t5 0.583833
R317 a_5381_1389.n1 a_5381_1389.t11 0.583833
R318 a_5381_1389.n0 a_5381_1389.t16 0.583833
R319 a_5381_1389.n0 a_5381_1389.t19 0.583833
R320 a_5381_1389.n17 a_5381_1389.t9 0.583833
R321 a_5381_1389.t18 a_5381_1389.n17 0.583833
R322 a_5381_1389.n4 a_5381_1389.n2 0.06818
R323 a_5381_1389.n6 a_5381_1389.n4 0.06818
R324 a_5381_1389.n8 a_5381_1389.n6 0.06818
R325 a_5381_1389.n10 a_5381_1389.n8 0.06818
R326 a_5381_1389.n12 a_5381_1389.n10 0.06818
R327 a_5381_1389.n14 a_5381_1389.n12 0.06818
R328 a_5381_1389.n16 a_5381_1389.n14 0.06818
R329 vdd.t1 vdd.t24 1159.16
R330 vdd.t2 vdd.t26 1138.89
R331 vdd.t23 vdd.t31 1132.35
R332 vdd.t29 vdd.n9 888.654
R333 vdd.n2 vdd.t23 522.399
R334 vdd.n10 vdd.t29 522.338
R335 vdd.t24 vdd.n0 522.337
R336 vdd.t31 vdd.n1 517.273
R337 vdd.n1 vdd.t0 517.273
R338 vdd.t26 vdd.n8 517.273
R339 vdd.n8 vdd.t1 517.273
R340 vdd.n9 vdd.t2 513.072
R341 vdd.n4 vdd.t19 304.387
R342 vdd.t19 vdd.t22 208.889
R343 vdd.t22 vdd.t8 208.889
R344 vdd.t8 vdd.t14 208.889
R345 vdd.t14 vdd.t4 208.889
R346 vdd.t4 vdd.t15 208.889
R347 vdd.t15 vdd.t20 208.889
R348 vdd.t20 vdd.t7 208.889
R349 vdd.t7 vdd.t10 208.889
R350 vdd.t10 vdd.t17 208.889
R351 vdd.t17 vdd.t11 208.889
R352 vdd.t11 vdd.t18 208.889
R353 vdd.t18 vdd.t5 208.889
R354 vdd.t5 vdd.t9 208.889
R355 vdd.t9 vdd.t16 208.889
R356 vdd.t16 vdd.t3 208.889
R357 vdd.t3 vdd.t12 208.889
R358 vdd.t12 vdd.t21 208.889
R359 vdd.t21 vdd.t6 208.889
R360 vdd.t6 vdd.t13 208.889
R361 vdd.n6 vdd.t28 9.66464
R362 vdd.n14 vdd.n0 7.11612
R363 vdd.n9 vdd.n5 6.96188
R364 vdd.n2 vdd.n1 6.29206
R365 vdd.n0 vdd.t25 5.262
R366 vdd.n10 vdd.t30 5.26126
R367 vdd.n6 vdd.t27 3.69646
R368 vdd.n4 vdd.n3 3.54271
R369 vdd.n8 vdd.n7 3.13374
R370 vdd.n11 vdd.n10 2.43993
R371 vdd.n13 vdd.n3 2.17281
R372 vdd.n12 vdd.n4 2.08974
R373 vdd.n14 vdd.n13 1.68062
R374 vdd.n7 vdd.n6 1.60498
R375 vdd.n3 vdd.n2 0.698
R376 vdd.n7 vdd.n5 0.337689
R377 vdd.n11 vdd.n5 0.248933
R378 vdd.n13 vdd.n12 0.206214
R379 vdd vdd.n14 0.157631
R380 vdd.n12 vdd.n11 0.0067212
R381 clk.n3 clk.t0 35.7254
R382 clk.n0 clk.t6 35.7221
R383 clk.n5 clk.t5 34.1136
R384 clk.n4 clk.t1 30.1393
R385 clk.n1 clk.t4 30.1393
R386 clk.n2 clk.t2 27.1236
R387 clk.n3 clk.t3 15.823
R388 clk.n0 clk.t7 15.8225
R389 clk.n1 clk.n0 10.6732
R390 clk.n4 clk.n3 10.6727
R391 clk.n6 clk.n2 1.52712
R392 clk clk.n6 0.460065
R393 clk.n6 clk.n5 0.281711
R394 clk.n2 clk.n1 0.111676
R395 clk.n5 clk.n4 0.0995311
R396 vin.n0 vin.t3 13.8016
R397 vin.n7 vin.t2 9.92542
R398 vin vin.n6 9.75035
R399 vin.n1 vin.n0 4.99212
R400 vin.n3 vin.n2 4.60986
R401 vin.n4 vin.n3 4.5696
R402 vin.n5 vin.n4 4.5005
R403 vin.n2 vin.n1 4.5005
R404 vin.n3 vin.t0 3.48383
R405 vin.n7 vin.t1 3.48383
R406 vin.n6 vin.n5 1.04563
R407 vin.n6 vin 0.722519
R408 vin vin.n7 0.394842
R409 vin.n5 vin.n1 0.1805
R410 vin.n4 vin 0.096125
R411 vin.n2 vin 0.084875
R412 vin.n0 vin 0.037625
R413 nclk.n0 nclk.t7 35.0711
R414 nclk.n3 nclk.t1 28.37
R415 nclk.n1 nclk.t6 25.9811
R416 nclk.n3 nclk.t0 25.2836
R417 nclk.n5 nclk.t4 24.2876
R418 nclk.n2 nclk.t3 24.2876
R419 nclk.n4 nclk.t2 19.9399
R420 nclk.n0 nclk.t5 19.5588
R421 nclk.n2 nclk.n1 7.06888
R422 nclk.n5 nclk.n4 7.0647
R423 nclk.n6 nclk.n5 2.40549
R424 nclk.n6 nclk.n2 1.7803
R425 nclk.n4 nclk.n3 0.699125
R426 nclk nclk.n6 0.594832
R427 nclk.n1 nclk.n0 0.381269
C0 a_8034_n1134# a_5673_n171# 0.31123f
C1 vout vdd 1.94401f
C2 a_5944_2887# vdd 0.3862f
C3 vin vout 2.42574f
C4 a_5673_n171# vdd 1.3089f
C5 clk vout 1.05144f
C6 a_8034_n1134# vdd 0.5497f
C7 a_8039_2775# vout 0.00196f
C8 vin a_5944_2887# 0.05549f
C9 a_5944_2887# clk 0.87934f
C10 a_5944_2887# a_8039_2775# 0.87223f
C11 vin a_5673_n171# 0.43115f
C12 vin a_8034_n1134# 0.23324f
C13 clk a_5673_n171# 0.74034f
C14 clk a_8034_n1134# 0.65791f
C15 nclk vout 0.17473f
C16 a_5944_2887# nclk 0.12006f
C17 vin vdd 1.17738f
C18 clk vdd 2.16069f
C19 nclk a_5673_n171# 0.93861f
C20 a_8039_2775# vdd 0.86692f
C21 a_8034_n1134# nclk 0.5632f
C22 vin clk 0.13047f
C23 vin a_8039_2775# 0.50625f
C24 a_5904_n1280# vout 0.00174f
C25 clk a_8039_2775# 0.68185f
C26 a_5904_n1280# a_5673_n171# 0.78751f
C27 a_8034_n1134# a_5904_n1280# 0.91362f
C28 nclk vdd 3.21794f
C29 vin nclk 0.69675f
C30 clk nclk 2.7322f
C31 nclk a_8039_2775# 0.68724f
C32 a_5904_n1280# vdd 0.23322f
C33 vin a_5904_n1280# 0.02438f
C34 clk a_5904_n1280# 0.82417f
C35 a_5904_n1280# nclk 0.12185f
C36 a_5944_2887# vout 0.00216f
C37 a_5673_n171# vout 1.37316f
C38 a_8034_n1134# vout 0.00218f
C39 vout vss 5.0405f
C40 vin vss 3.03134f
C41 nclk vss 6.76573f
C42 clk vss 8.65105f
C43 vdd vss 41.01737f
C44 a_8034_n1134# vss 4.47584f
C45 a_5904_n1280# vss 2.55107f
C46 a_5673_n171# vss 4.27103f
C47 a_8039_2775# vss 2.74755f
C48 a_5944_2887# vss 1.5224f
C49 nclk.t7 vss 0.02839f
C50 nclk.t5 vss 0.1214f
C51 nclk.n0 vss 0.25404f
C52 nclk.t6 vss 0.13476f
C53 nclk.n1 vss 0.48461f
C54 nclk.t3 vss 0.16661f
C55 nclk.n2 vss 0.58828f
C56 nclk.t2 vss 0.12284f
C57 nclk.t1 vss 0.02302f
C58 nclk.t0 vss 0.12928f
C59 nclk.n3 vss 0.48242f
C60 nclk.n4 vss 0.35941f
C61 nclk.t4 vss 0.16661f
C62 nclk.n5 vss 0.7867f
C63 nclk.n6 vss 1.61769f
C64 vin.t3 vss 0.02556f
C65 vin.n0 vss 0.01809f
C66 vin.n1 vss 0.0555f
C67 vin.n2 vss 0.00832f
C68 vin.t0 vss 0.03762f
C69 vin.n3 vss 0.04102f
C70 vin.n4 vss 0.00868f
C71 vin.n5 vss 0.05685f
C72 vin.n6 vss 6.55048f
C73 vin.t2 vss 0.02324f
C74 vin.t1 vss 0.03762f
C75 vin.n7 vss 0.09641f
C76 clk.t2 vss 0.00995f
C77 clk.t7 vss 0.04631f
C78 clk.t6 vss 0.12799f
C79 clk.n0 vss 0.30308f
C80 clk.t4 vss 0.14359f
C81 clk.n1 vss 0.45504f
C82 clk.n2 vss 0.91656f
C83 clk.t5 vss 0.01691f
C84 clk.t3 vss 0.04631f
C85 clk.t0 vss 0.13424f
C86 clk.n3 vss 0.30815f
C87 clk.t1 vss 0.14359f
C88 clk.n4 vss 0.4463f
C89 clk.n5 vss 0.29462f
C90 clk.n6 vss 1.13327f
C91 vdd.t25 vss 0.01441f
C92 vdd.n0 vss 0.15444f
C93 vdd.t0 vss 0.23274f
C94 vdd.n1 vss 0.43568f
C95 vdd.t31 vss 0.23024f
C96 vdd.t23 vss 0.2318f
C97 vdd.n2 vss 0.23013f
C98 vdd.n3 vss -0.16687f
C99 vdd.t13 vss 0.27036f
C100 vdd.t6 vss 0.12581f
C101 vdd.t21 vss 0.12581f
C102 vdd.t12 vss 0.12581f
C103 vdd.t3 vss 0.12581f
C104 vdd.t16 vss 0.12581f
C105 vdd.t9 vss 0.12581f
C106 vdd.t5 vss 0.12581f
C107 vdd.t18 vss 0.12581f
C108 vdd.t11 vss 0.12581f
C109 vdd.t17 vss 0.12581f
C110 vdd.t10 vss 0.12581f
C111 vdd.t7 vss 0.12581f
C112 vdd.t20 vss 0.12581f
C113 vdd.t15 vss 0.12581f
C114 vdd.t4 vss 0.12581f
C115 vdd.t14 vss 0.12581f
C116 vdd.t8 vss 0.12581f
C117 vdd.t22 vss 0.12581f
C118 vdd.t19 vss 0.1552f
C119 vdd.n4 vss 0.25697f
C120 vdd.n5 vss 0.13103f
C121 vdd.t24 vss 0.17018f
C122 vdd.t1 vss 0.22035f
C123 vdd.t28 vss 0.01263f
C124 vdd.t27 vss 0.0231f
C125 vdd.n6 vss 0.06737f
C126 vdd.n7 vss 0.12697f
C127 vdd.n8 vss 0.43367f
C128 vdd.t26 vss 0.23115f
C129 vdd.t2 vss 0.23003f
C130 vdd.n9 vss 0.16748f
C131 vdd.t29 vss 0.13653f
C132 vdd.t30 vss 0.01444f
C133 vdd.n10 vss 0.13085f
C134 vdd.n11 vss 0.09682f
C135 vdd.n12 vss 0.08416f
C136 vdd.n13 vss 1.5051f
C137 vdd.n14 vss 1.1739f
C138 a_5381_1389.t9 vss 0.06811f
C139 a_5381_1389.t16 vss 0.06811f
C140 a_5381_1389.t19 vss 0.06811f
C141 a_5381_1389.n0 vss 0.2315f
C142 a_5381_1389.t5 vss 0.06811f
C143 a_5381_1389.t11 vss 0.06811f
C144 a_5381_1389.n1 vss 0.21423f
C145 a_5381_1389.n2 vss 1.37545f
C146 a_5381_1389.t1 vss 0.06811f
C147 a_5381_1389.t12 vss 0.06811f
C148 a_5381_1389.n3 vss 0.21423f
C149 a_5381_1389.n4 vss 0.85169f
C150 a_5381_1389.t17 vss 0.06811f
C151 a_5381_1389.t4 vss 0.06811f
C152 a_5381_1389.n5 vss 0.21423f
C153 a_5381_1389.n6 vss 0.85169f
C154 a_5381_1389.t7 vss 0.06811f
C155 a_5381_1389.t14 vss 0.06811f
C156 a_5381_1389.n7 vss 0.21423f
C157 a_5381_1389.n8 vss 0.85169f
C158 a_5381_1389.t8 vss 0.06811f
C159 a_5381_1389.t15 vss 0.06811f
C160 a_5381_1389.n9 vss 0.21423f
C161 a_5381_1389.n10 vss 0.85169f
C162 a_5381_1389.t2 vss 0.06811f
C163 a_5381_1389.t6 vss 0.06811f
C164 a_5381_1389.n11 vss 0.21423f
C165 a_5381_1389.n12 vss 0.85169f
C166 a_5381_1389.t13 vss 0.06811f
C167 a_5381_1389.t0 vss 0.06811f
C168 a_5381_1389.n13 vss 0.21423f
C169 a_5381_1389.n14 vss 0.85169f
C170 a_5381_1389.t3 vss 0.06811f
C171 a_5381_1389.t10 vss 0.06811f
C172 a_5381_1389.n15 vss 0.2315f
C173 a_5381_1389.n16 vss 1.37546f
C174 a_5381_1389.n17 vss 0.21422f
C175 a_5381_1389.t18 vss 0.06811f
C176 a_5297_1329.t1 vss 0.06065f
C177 a_5297_1329.n2 vss 0.02076f
C178 a_5297_1329.t13 vss 0.0822f
C179 a_5297_1329.t20 vss 0.08194f
C180 a_5297_1329.n3 vss 0.11187f
C181 a_5297_1329.t5 vss 0.08194f
C182 a_5297_1329.n4 vss 0.06021f
C183 a_5297_1329.t14 vss 0.08194f
C184 a_5297_1329.n5 vss 0.06021f
C185 a_5297_1329.t23 vss 0.08194f
C186 a_5297_1329.n6 vss 0.06021f
C187 a_5297_1329.t10 vss 0.08194f
C188 a_5297_1329.n7 vss 0.06021f
C189 a_5297_1329.t17 vss 0.08194f
C190 a_5297_1329.n8 vss 0.06021f
C191 a_5297_1329.t21 vss 0.08194f
C192 a_5297_1329.n9 vss 0.05331f
C193 a_5297_1329.n10 vss 0.02078f
C194 a_5297_1329.t15 vss 0.08194f
C195 a_5297_1329.n11 vss 0.04715f
C196 a_5297_1329.t8 vss 0.08194f
C197 a_5297_1329.n12 vss 0.04714f
C198 a_5297_1329.n13 vss 0.02078f
C199 a_5297_1329.t7 vss 0.0822f
C200 a_5297_1329.t4 vss 0.08194f
C201 a_5297_1329.n14 vss 0.11187f
C202 a_5297_1329.t18 vss 0.08194f
C203 a_5297_1329.n15 vss 0.06021f
C204 a_5297_1329.t12 vss 0.08194f
C205 a_5297_1329.n16 vss 0.06021f
C206 a_5297_1329.t22 vss 0.08194f
C207 a_5297_1329.n17 vss 0.06021f
C208 a_5297_1329.t11 vss 0.08194f
C209 a_5297_1329.n18 vss 0.06021f
C210 a_5297_1329.t6 vss 0.08194f
C211 a_5297_1329.n19 vss 0.06021f
C212 a_5297_1329.t19 vss 0.08194f
C213 a_5297_1329.n20 vss 0.06021f
C214 a_5297_1329.t16 vss 0.08194f
C215 a_5297_1329.n21 vss 0.05059f
C216 a_5297_1329.t9 vss 0.08194f
C217 a_5297_1329.n22 vss 0.04717f
C218 a_5297_1329.n23 vss 0.02074f
C219 a_5297_1329.n24 vss 0.76429f
C220 a_5297_1329.n25 vss 0.19448f
C221 a_5297_1329.t2 vss 0.06065f
C222 a_5297_1329.t3 vss 0.03285f
C223 a_5297_1329.n26 vss 0.14217f
C224 a_5297_1329.n27 vss 0.36174f
C225 a_5297_1329.n28 vss 0.19448f
C226 a_5297_1329.n29 vss 0.17367f
C227 a_5297_1329.n30 vss 0.82621f
C228 a_5297_1329.n31 vss 0.16023f
C229 a_5297_1329.n32 vss 0.14199f
C230 a_5297_1329.t0 vss 0.03285f
C231 vout.n0 vss 0.11453f
C232 vout.t21 vss 0.27416f
C233 vout.t5 vss 0.22981f
C234 vout.n1 vss 0.71753f
C235 vout.t24 vss 0.04819f
C236 vout.t29 vss 0.04819f
C237 vout.n2 vss 0.1478f
C238 vout.t1 vss 0.04819f
C239 vout.t4 vss 0.04819f
C240 vout.n3 vss 0.1478f
C241 vout.t6 vss 0.06047f
C242 vout.t11 vss 0.06047f
C243 vout.n4 vss 0.18419f
C244 vout.n5 vss 0.33623f
C245 vout.n6 vss 0.11453f
C246 vout.t0 vss 0.04819f
C247 vout.t2 vss 0.04819f
C248 vout.n7 vss 0.1478f
C249 vout.t14 vss 0.06047f
C250 vout.t18 vss 0.06047f
C251 vout.n8 vss 0.18419f
C252 vout.n9 vss 0.11405f
C253 vout.n10 vss 0.11453f
C254 vout.t28 vss 0.04819f
C255 vout.t25 vss 0.04819f
C256 vout.n11 vss 0.1478f
C257 vout.t7 vss 0.06047f
C258 vout.t10 vss 0.06047f
C259 vout.n12 vss 0.18419f
C260 vout.t3 vss 0.04819f
C261 vout.t27 vss 0.04819f
C262 vout.n13 vss 0.1478f
C263 vout.t15 vss 0.06047f
C264 vout.t16 vss 0.06047f
C265 vout.n14 vss 0.18419f
C266 vout.n15 vss 0.33623f
C267 vout.n16 vss 0.11453f
C268 vout.t22 vss 0.04819f
C269 vout.t23 vss 0.04819f
C270 vout.n17 vss 0.1478f
C271 vout.t19 vss 0.06047f
C272 vout.t9 vss 0.06047f
C273 vout.n18 vss 0.18419f
C274 vout.n19 vss 0.11405f
C275 vout.n20 vss 0.11453f
C276 vout.t33 vss 0.04819f
C277 vout.t35 vss 0.04819f
C278 vout.n21 vss 0.1478f
C279 vout.t12 vss 0.06047f
C280 vout.t17 vss 0.06047f
C281 vout.n22 vss 0.18419f
C282 vout.t34 vss 0.04819f
C283 vout.t26 vss 0.04819f
C284 vout.n23 vss 0.1478f
C285 vout.t20 vss 0.06047f
C286 vout.t8 vss 0.06047f
C287 vout.n24 vss 0.18419f
C288 vout.n25 vss 0.33623f
C289 vout.n26 vss 0.20378f
C290 vout.t32 vss 0.04819f
C291 vout.t31 vss 0.04819f
C292 vout.n27 vss 0.1478f
C293 vout.t13 vss 0.27416f
C294 vout.t30 vss 0.22981f
C295 vout.n28 vss 0.7161f
C296 vout.n29 vss 0.01235f
C297 vout.n30 vss 0.18821f
C298 vout.n31 vss 0.10764f
C299 vout.n32 vss 0.0834f
C300 vout.n33 vss 0.11453f
C301 vout.n34 vss 0.11453f
C302 vout.n35 vss 0.08768f
C303 vout.n36 vss 0.10336f
C304 vout.n37 vss 0.33623f
C305 vout.n38 vss 0.06772f
C306 vout.n39 vss 0.11453f
C307 vout.n40 vss 0.11453f
C308 vout.n41 vss 0.11453f
C309 vout.n42 vss 0.06629f
C310 vout.n43 vss 0.33623f
C311 vout.n44 vss 0.10479f
C312 vout.n45 vss 0.08625f
C313 vout.n46 vss 0.11453f
C314 vout.n47 vss 0.11453f
C315 vout.n48 vss 0.08483f
C316 vout.n49 vss 0.10621f
C317 vout.n50 vss 0.33623f
C318 vout.n51 vss 0.06487f
C319 vout.n52 vss 0.11453f
C320 vout.n53 vss 0.11453f
C321 vout.n54 vss 0.11453f
C322 vout.n55 vss 0.06914f
C323 vout.n56 vss 0.33623f
C324 vout.n57 vss 0.10193f
C325 vout.n58 vss 0.0891f
C326 vout.n59 vss 0.11453f
C327 vout.n60 vss 0.11453f
C328 vout.n61 vss 0.08197f
C329 vout.n62 vss 0.10906f
C330 vout.n63 vss 0.18821f
C331 vout.n64 vss 0.00998f
C332 vout.n65 vss 1.03825f
C333 a_5757_n39.t11 vss 0.06767f
C334 a_5757_n39.t5 vss 0.06767f
C335 a_5757_n39.t3 vss 0.06767f
C336 a_5757_n39.n0 vss 0.22789f
C337 a_5757_n39.t7 vss 0.06767f
C338 a_5757_n39.t10 vss 0.06767f
C339 a_5757_n39.n1 vss 0.22789f
C340 a_5757_n39.t14 vss 0.06767f
C341 a_5757_n39.t4 vss 0.06767f
C342 a_5757_n39.n2 vss 0.21228f
C343 a_5757_n39.n3 vss 1.43169f
C344 a_5757_n39.t8 vss 0.06767f
C345 a_5757_n39.t1 vss 0.06767f
C346 a_5757_n39.n4 vss 0.21228f
C347 a_5757_n39.n5 vss 0.88109f
C348 a_5757_n39.t13 vss 0.06767f
C349 a_5757_n39.t2 vss 0.06767f
C350 a_5757_n39.n6 vss 0.21228f
C351 a_5757_n39.n7 vss 0.88109f
C352 a_5757_n39.t9 vss 0.06767f
C353 a_5757_n39.t12 vss 0.06767f
C354 a_5757_n39.n8 vss 0.21228f
C355 a_5757_n39.n9 vss 0.88109f
C356 a_5757_n39.t15 vss 0.06767f
C357 a_5757_n39.t6 vss 0.06767f
C358 a_5757_n39.n10 vss 0.21228f
C359 a_5757_n39.n11 vss 0.88109f
C360 a_5757_n39.n12 vss 1.4317f
C361 a_5757_n39.n13 vss 0.21227f
C362 a_5757_n39.t0 vss 0.06767f
.ends

