magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l33d0 >>
<< l34d0 >>
<< l30d0 >>
<< l22d0 >>
<< l31d0 >>
<< l21d0 >>
<< labels >>
rlabel l34d10 -0.096 0.061 -0.096 0.061 0 
<< end >>
