* NGSPICE file created from swmatrix_row_10.ext - technology: gf180mcuD
.subckt swmatrix_row_10_pex D_out D_in PHI_1 PHI_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] VDD
+ pin VSS
X0 BUS[5].t16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 pin.t25 vdd.t88 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1 swmatrix_Tgate_3.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t428 vdd.t427 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X2 vdd.t71 a_51256_2002# a_51116_2122# vdd.t70 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X3 a_26296_2002# a_25952_2122# vss.t307 vss.t306 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X4 a_34508_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t289 vss.t288 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X5 BUS[8].t7 swmatrix_Tgate_3.gated_control pin.t15 vss.t22 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X6 a_53620_1577# a_52392_1562# a_53376_2122# vss.t206 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X7 pin.t194 swmatrix_Tgate_9.gated_control BUS[1].t17 vss.t342 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X8 a_6716_1580# a_6248_1562# vss.t250 vss.t249 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X9 pin.t52 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 BUS[3].t22 vdd.t113 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X10 BUS[1].t8 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 pin.t88 vdd.t228 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X11 vdd.t146 phi_2.t0 a_39912_1562# vdd.t145 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X12 pin.t229 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 BUS[8].t22 vdd.t525 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X13 pin.t212 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 BUS[6].t16 vdd.t493 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X14 a_4921_1539# ShiftReg_row_10_2$1_0.Q[1] vss.t330 vss.t329 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X15 vdd.t151 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t150 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X16 pin.t46 swmatrix_Tgate_2.gated_control BUS[10].t5 vss.t74 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X17 vss.t188 a_45016_2002# a_44916_1577# vss.t187 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X18 vdd.t272 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] vdd.t271 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X19 vss.t252 a_38776_2002# a_38676_1577# vss.t251 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X20 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t0 a_11161_1539# vss.t13 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X21 BUS[8].t0 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 pin.t6 vdd.t13 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X22 a_44156_1580# a_43688_1562# vss.t110 vss.t109 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X23 a_13472_2122# a_12488_1562# a_13324_2122# vdd.t61 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X24 a_19564_2122# ShiftReg_row_10_2$1_0.Q[3] vdd.t512 vdd.t511 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X25 vdd.t58 a_53720_2002# a_53580_2122# vdd.t57 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X26 BUS[2].t16 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 pin.t220 vdd.t507 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X27 vss.t315 phi_1.t0 a_56168_1562# vss.t314 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X28 vdd.t22 enable.t1 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t21 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X29 a_26156_2122# a_25436_1580# a_25952_2122# vdd.t391 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X30 a_56636_1580# a_56168_1562# vdd.t475 vdd.t474 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X31 a_19916_2122# a_19196_1580# a_19712_2122# vdd.t110 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X32 swmatrix_Tgate_7.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t112 vdd.t111 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X33 pin.t159 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 BUS[4].t16 vdd.t356 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X34 BUS[1].t5 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 pin.t85 vdd.t225 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X35 pin.t77 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 BUS[2].t15 vdd.t195 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X36 vdd.t495 phi_1.t1 a_12488_1562# vdd.t494 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X37 a_7576_2002# a_7232_2122# vdd.t241 vdd.t240 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X38 swmatrix_Tgate_2.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t411 vdd.t410 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X39 swmatrix_Tgate_1.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t141 vss.t140 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X40 vss.t220 a_47480_2002# a_47380_1577# vss.t219 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X41 vdd.t497 phi_1.t2 a_8_1562# vdd.t496 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X42 vss.t73 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t72 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X43 pin.t86 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[1].t6 vdd.t226 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X44 a_48601_1539# ShiftReg_row_10_2$1_0.Q[8] vss.t322 vss.t321 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X45 a_46620_1580# a_46152_1562# vss.t318 vss.t317 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X46 BUS[6].t15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 pin.t152 vdd.t349 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X47 vss.t105 phi_2.t1 a_58632_1562# vss.t104 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X48 a_34900_1577# a_33672_1562# a_34656_2122# vss.t158 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X49 a_28620_2122# a_27900_1580# a_28416_2122# vdd.t62 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X50 pin.t53 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 BUS[3].t21 vdd.t114 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X51 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[5] vdd.t157 vdd.t156 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X52 vss.t256 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t255 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X53 pin.t147 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 BUS[10].t16 vdd.t327 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X54 vss.t305 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t304 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X55 pin.t7 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[8].t1 vdd.t14 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X56 pin.t142 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 BUS[4].t15 vdd.t322 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X57 a_45016_2002# a_44672_2122# vdd.t18 vdd.t17 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X58 vss.t384 phi_1.t3 a_8_1562# vss.t383 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X59 pin.t209 swmatrix_Tgate_1.gated_control BUS[9].t21 vss.t380 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X60 vdd.t380 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t379 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X61 vss.t107 phi_2.t2 a_2472_1562# vss.t106 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X62 vdd.t31 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t30 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X63 a_32044_2122# ShiftReg_row_10_2$1_0.Q[5] vdd.t155 vdd.t154 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X64 BUS[10].t6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 pin.t80 vdd.t213 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X65 vss.t126 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t125 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X66 a_2940_1580# a_2472_1562# vdd.t99 vdd.t98 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X67 BUS[8].t16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 pin.t113 vdd.t281 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X68 a_53376_2122# a_52860_1580# a_53228_1577# vss.t290 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X69 BUS[4].t14 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 pin.t143 vdd.t323 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X70 BUS[9].t8 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 pin.t148 vdd.t339 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X71 BUS[7].t16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 pin.t165 vdd.t366 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X72 vdd.t199 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t198 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X73 swmatrix_Tgate_5.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t85 vss.t84 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X74 BUS[3].t5 swmatrix_Tgate_4.gated_control pin.t174 vss.t264 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X75 a_28760_2002# a_28416_2122# vss.t247 vss.t246 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X76 pin.t153 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[6].t14 vdd.t350 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X77 pin.t0 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[2].t14 vdd.t0 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X78 BUS[1].t7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 pin.t87 vdd.t227 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X79 a_47480_2002# a_47136_2122# vdd.t207 vdd.t206 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X80 vss.t359 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] vss.t358 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X81 a_23641_1539# ShiftReg_row_10_2$1_0.Q[4] vss.t199 vss.t198 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X82 vss.t235 phi_2.t3 a_39912_1562# vss.t234 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X83 pin.t124 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 BUS[9].t4 vdd.t298 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X84 a_7084_1577# ShiftReg_row_10_2$1_0.Q[1] vss.t328 vss.t327 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X85 a_1336_2002# a_992_2122# vss.t89 vss.t88 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X86 vdd.t56 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] vdd.t55 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X87 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[2] vdd.t41 vdd.t40 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X88 vdd.t124 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] vdd.t123 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X89 BUS[2].t13 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 pin.t1 vdd.t1 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X90 a_61081_1539# d_out.t2 vss.t233 vss.t232 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X91 pin.t60 swmatrix_Tgate_5.gated_control BUS[5].t22 vss.t118 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X92 BUS[8].t17 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t114 vdd.t282 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X93 a_27900_1580# a_27432_1562# vss.t92 vss.t91 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X94 BUS[5].t15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 pin.t31 vdd.t87 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X95 vss.t379 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t378 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X96 BUS[3].t20 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 pin.t19 vdd.t45 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X97 vdd.t219 a_59616_2122# d_out.t1 vdd.t218 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X98 a_32192_2122# a_31676_1580# a_32044_1577# vss.t231 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X99 a_25952_2122# a_25436_1580# a_25804_1577# vss.t275 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X100 BUS[7].t22 swmatrix_Tgate_0.gated_control pin.t217 vss.t392 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X101 pin.t81 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[10].t7 vdd.t214 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X102 a_44524_1577# ShiftReg_row_10_2$1_0.Q[7] vss.t274 vss.t273 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X103 pin.t199 swmatrix_Tgate_9.gated_control BUS[1].t16 vss.t341 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X104 vdd.t445 phi_1.t4 a_49928_1562# vdd.t444 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X105 vdd.t462 enable.t2 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t461 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X106 pin.t27 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[5].t14 vdd.t86 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X107 vdd.t464 enable.t3 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t463 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X108 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t4 a_48601_1539# vss.t345 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X109 vss.t324 phi_1.t5 a_12488_1562# vss.t323 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X110 pin.t125 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 BUS[9].t5 vdd.t299 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X111 a_59468_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t501 vdd.t500 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X112 a_53376_2122# a_52392_1562# a_53228_2122# vdd.t280 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X113 pin.t216 swmatrix_Tgate_0.gated_control BUS[7].t21 vss.t391 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X114 a_12956_1580# a_12488_1562# vdd.t60 vdd.t59 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X115 a_22520_2002# a_22176_2122# vdd.t54 vdd.t53 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X116 pin.t14 swmatrix_Tgate_3.gated_control BUS[8].t6 vss.t21 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X117 BUS[9].t22 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 pin.t221 vdd.t508 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X118 a_45016_2002# a_44672_2122# vss.t10 vss.t9 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X119 vss.t117 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t116 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X120 a_46988_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t155 vss.t154 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X121 a_41240_2002# a_40896_2122# vss.t287 vss.t286 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X122 a_844_2122# D_in.t0 vdd.t517 vdd.t516 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X123 vss.t160 a_10040_2002# a_9940_1577# vss.t159 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X124 pin.t2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 BUS[2].t12 vdd.t2 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X125 BUS[10].t4 swmatrix_Tgate_2.gated_control pin.t45 vss.t71 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X126 vdd.t344 phi_2.t4 a_52392_1562# vdd.t343 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X127 vss.t237 phi_2.t5 a_21192_1562# vss.t236 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X128 vdd.t94 a_35000_2002# a_34860_2122# vdd.t93 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X129 swmatrix_Tgate_9.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t173 vdd.t172 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X130 pin.t26 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[5].t13 vdd.t85 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X131 pin.t20 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[3].t19 vdd.t46 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X132 a_21660_1580# a_21192_1562# vdd.t260 vdd.t259 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X133 pin.t189 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[10].t22 vdd.t422 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X134 pin.t44 swmatrix_Tgate_2.gated_control BUS[10].t3 vss.t70 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X135 vss.t174 a_57496_2002# a_57396_1577# vss.t173 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X136 a_38284_2122# ShiftReg_row_10_2$1_0.Q[6] vdd.t294 vdd.t293 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X137 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[1] vdd.t449 vdd.t448 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X138 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t5 a_23641_1539# vss.t11 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X139 a_32192_2122# a_31208_1562# a_32044_2122# vdd.t140 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X140 a_56636_1580# a_56168_1562# vss.t353 vss.t352 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X141 a_9180_1580# a_8712_1562# vdd.t421 vdd.t420 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X142 a_25952_2122# a_24968_1562# a_25804_2122# vdd.t418 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X143 BUS[5].t12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t40 vdd.t84 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X144 a_34508_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t402 vdd.t401 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X145 BUS[3].t18 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t21 vdd.t47 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X146 BUS[10].t19 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t162 vdd.t359 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X147 a_44916_1577# a_43688_1562# a_44672_2122# vss.t108 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X148 a_38636_2122# a_37916_1580# a_38432_2122# vdd.t169 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X149 BUS[2].t22 swmatrix_Tgate_8.gated_control pin.t67 vss.t124 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X150 BUS[2].t11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t3 vdd.t3 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X151 a_25804_1577# ShiftReg_row_10_2$1_0.Q[4] vss.t197 vss.t196 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X152 vss.t334 a_1336_2002# a_1236_1577# vss.t333 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X153 a_20056_2002# a_19712_2122# vss.t55 vss.t54 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X154 a_22028_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t144 vss.t143 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X155 pin.t154 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[6].t13 vdd.t351 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X156 a_16180_1577# a_14952_1562# a_15936_2122# vss.t223 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X157 pin.t130 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[4].t13 vdd.t310 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X158 pin.t69 swmatrix_Tgate_8.gated_control BUS[2].t21 vss.t123 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X159 a_9548_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t34 vss.t33 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X160 BUS[8].t18 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t115 vdd.t283 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X161 BUS[6].t12 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t22 vdd.t48 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X162 vss.t263 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t262 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X163 BUS[3].t17 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t89 vdd.t229 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X164 pin.t16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 BUS[1].t0 vdd.t42 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X165 a_47340_2122# a_46620_1580# a_47136_2122# vdd.t486 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X166 a_22520_2002# a_22176_2122# vss.t38 vss.t37 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X167 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[8] vdd.t443 vdd.t442 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X168 a_13324_2122# ShiftReg_row_10_2$1_0.Q[2] vdd.t39 vdd.t38 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X169 vss.t8 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t7 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X170 vss.t297 a_3800_2002# a_3700_1577# vss.t296 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X171 vdd.t346 phi_2.t6 a_33672_1562# vdd.t345 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X172 vss.t326 phi_1.t6 a_49928_1562# vss.t325 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X173 a_28416_2122# a_27900_1580# a_28268_1577# vss.t44 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X174 pin.t35 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 BUS[5].t11 vdd.t83 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X175 a_57496_2002# a_57152_2122# vdd.t103 vdd.t102 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X176 a_2940_1580# a_2472_1562# vss.t62 vss.t61 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X177 vdd.t135 a_16280_2002# a_16140_2122# vdd.t134 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X178 BUS[9].t20 swmatrix_Tgate_1.gated_control pin.t208 vss.t377 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X179 vdd.t378 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t377 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X180 vdd.t426 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t425 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X181 a_50764_2122# ShiftReg_row_10_2$1_0.Q[8] vdd.t441 vdd.t440 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X182 pin.t126 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 BUS[7].t15 vdd.t304 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X183 a_19196_1580# a_18728_1562# vdd.t160 vdd.t159 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X184 a_7476_1577# a_6248_1562# a_7232_2122# vss.t248 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X185 BUS[5].t10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 pin.t34 vdd.t82 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X186 a_37916_1580# a_37448_1562# vss.t228 vss.t227 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X187 pin.t211 swmatrix_Tgate_1.gated_control BUS[9].t19 vss.t376 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X188 a_15788_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t471 vdd.t470 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X189 a_1336_2002# a_992_2122# vdd.t130 vdd.t129 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X190 BUS[9].t0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t78 vdd.t202 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X191 BUS[6].t11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t23 vdd.t49 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X192 BUS[4].t12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 pin.t131 vdd.t311 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X193 swmatrix_Tgate_0.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t398 vss.t397 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X194 BUS[4].t22 swmatrix_Tgate_7.gated_control pin.t205 vss.t369 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X195 vss.t270 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] vss.t269 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X196 pin.t4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[2].t10 vdd.t4 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X197 a_42361_1539# ShiftReg_row_10_2$1_0.Q[7] vss.t272 vss.t271 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X198 swmatrix_Tgate_4.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t120 vdd.t119 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X199 BUS[5].t21 swmatrix_Tgate_5.gated_control pin.t59 vss.t115 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X200 pin.t104 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[8].t13 vdd.t261 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X201 pin.t24 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[6].t10 vdd.t50 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X202 vdd.t481 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] vdd.t480 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X203 vdd.t222 a_7576_2002# a_7436_2122# vdd.t221 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X204 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[4] vdd.t268 vdd.t267 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X205 BUS[1].t15 swmatrix_Tgate_9.gated_control pin.t198 vss.t340 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X206 a_9940_1577# a_8712_1562# a_9696_2122# vss.t303 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X207 pin.t215 swmatrix_Tgate_0.gated_control BUS[7].t20 vss.t390 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X208 BUS[10].t20 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t163 vdd.t360 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X209 pin.t61 swmatrix_Tgate_5.gated_control BUS[5].t20 vss.t114 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X210 vdd.t20 enable.t6 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t19 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X211 BUS[8].t14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t105 vdd.t262 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X212 vss.t186 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t185 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X213 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out.t3 vdd.t341 vdd.t340 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X214 a_44672_2122# a_44156_1580# a_44524_1577# vss.t45 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X215 vss.t396 a_20056_2002# a_19956_1577# vss.t395 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X216 a_28416_2122# a_27432_1562# a_28268_2122# vdd.t133 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X217 BUS[9].t1 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t79 vdd.t203 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X218 BUS[7].t14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 pin.t136 vdd.t316 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X219 vss.t372 a_13816_2002# a_13716_1577# vss.t371 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X220 BUS[7].t19 swmatrix_Tgate_0.gated_control pin.t214 vss.t389 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X221 a_12956_1580# a_12488_1562# vss.t43 vss.t42 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X222 vss.t409 phi_1.t7 a_31208_1562# vss.t408 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X223 vdd.t251 a_45016_2002# a_44876_2122# vdd.t250 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X224 a_28268_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t172 vss.t171 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X225 a_38776_2002# a_38432_2122# vdd.t166 vdd.t165 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X226 pin.t187 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[9].t14 vdd.t414 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X227 a_31676_1580# a_31208_1562# vdd.t139 vdd.t138 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X228 pin.t137 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 BUS[7].t13 vdd.t317 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X229 a_41240_2002# a_40896_2122# vdd.t400 vdd.t399 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X230 BUS[2].t9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t5 vdd.t5 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X231 a_57496_2002# a_57152_2122# vss.t66 vss.t65 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X232 a_59960_2002# a_59616_2122# vss.t180 vss.t179 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X233 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t7 a_4921_1539# vss.t12 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X234 vss.t135 a_22520_2002# a_22420_1577# vss.t134 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X235 BUS[3].t16 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 pin.t90 vdd.t230 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X236 BUS[10].t17 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 pin.t157 vdd.t354 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X237 a_21660_1580# a_21192_1562# vss.t195 vss.t194 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X238 vss.t190 phi_2.t7 a_33672_1562# vss.t189 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X239 a_40380_1580# a_39912_1562# vdd.t406 vdd.t405 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X240 a_9180_1580# a_8712_1562# vss.t302 vss.t301 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X241 a_26196_1577# a_24968_1562# a_25952_2122# vss.t300 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X242 pin.t91 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 BUS[3].t15 vdd.t231 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X243 a_19956_1577# a_18728_1562# a_19712_2122# vss.t133 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X244 pin.t109 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 BUS[7].t12 vdd.t274 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X245 pin.t158 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 BUS[10].t18 vdd.t355 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X246 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t8 a_42361_1539# vss.t354 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X247 a_7232_2122# a_6716_1580# a_7084_1577# vss.t95 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X248 a_20056_2002# a_19712_2122# vdd.t92 vdd.t91 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X249 pin.t56 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[2].t8 vdd.t117 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X250 a_53228_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t201 vdd.t200 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X251 a_44672_2122# a_43688_1562# a_44524_2122# vdd.t149 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X252 vdd.t477 enable.t9 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t476 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X253 pin.t180 swmatrix_Tgate_6.gated_control BUS[6].t22 vss.t283 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X254 BUS[9].t15 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t188 vdd.t415 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X255 pin.t204 swmatrix_Tgate_7.gated_control BUS[4].t21 vss.t368 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X256 a_57356_2122# a_56636_1580# a_57152_2122# vdd.t472 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X257 BUS[7].t11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t110 vdd.t275 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X258 swmatrix_Tgate_1.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t168 vdd.t167 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X259 swmatrix_Tgate_3.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t309 vss.t308 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X260 BUS[4].t11 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t140 vdd.t320 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X261 a_3800_2002# a_3456_2122# vdd.t270 vdd.t269 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X262 a_32536_2002# a_32192_2122# vss.t254 vss.t253 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X263 a_40748_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t152 vss.t151 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X264 vdd.t527 phi_1.t8 a_43688_1562# vdd.t526 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X265 BUS[8].t5 swmatrix_Tgate_3.gated_control pin.t13 vss.t20 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X266 vdd.t455 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t454 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X267 BUS[6].t21 swmatrix_Tgate_6.gated_control pin.t179 vss.t282 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X268 vdd.t492 a_26296_2002# a_26156_2122# vdd.t491 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X269 a_9696_2122# a_9180_1580# a_9548_1577# vss.t175 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X270 a_28660_1577# a_27432_1562# a_28416_2122# vss.t90 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X271 pin.t190 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[3].t14 vdd.t430 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X272 a_59100_1580# a_58632_1562# vdd.t434 vdd.t433 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X273 BUS[1].t1 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 pin.t17 vdd.t43 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X274 a_1196_2122# a_476_1580# a_992_2122# vdd.t465 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X275 vss.t150 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] vss.t149 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X276 vdd.t253 phi_2.t8 a_14952_1562# vdd.t252 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X277 a_476_1580# a_8_1562# vdd.t8 vdd.t7 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X278 BUS[5].t9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t38 vdd.t81 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X279 pin.t210 swmatrix_Tgate_1.gated_control BUS[9].t18 vss.t375 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X280 BUS[3].t13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 pin.t191 vdd.t431 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X281 a_59820_2122# a_59100_1580# a_59616_2122# vdd.t456 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X282 pin.t18 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[1].t2 vdd.t44 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X283 BUS[8].t15 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 pin.t106 vdd.t263 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X284 a_25804_2122# ShiftReg_row_10_2$1_0.Q[4] vdd.t266 vdd.t265 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X285 a_47136_2122# a_46620_1580# a_46988_1577# vss.t370 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X286 BUS[2].t7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 pin.t57 vdd.t118 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X287 a_19196_1580# a_18728_1562# vss.t132 vss.t131 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X288 vdd.t96 a_28760_2002# a_28620_2122# vdd.t95 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X289 a_7232_2122# a_6248_1562# a_7084_2122# vdd.t370 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X290 vdd.t16 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t15 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X291 a_3660_2122# a_2940_1580# a_3456_2122# vdd.t215 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X292 pin.t54 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 BUS[8].t8 vdd.t115 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X293 pin.t192 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 BUS[4].t10 vdd.t438 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X294 vdd.t499 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t498 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X295 pin.t42 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[2].t6 vdd.t104 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X296 vss.t87 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t86 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X297 vss.t407 a_59960_2002# a_59860_1577# vss.t406 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X298 vdd.t529 phi_1.t9 a_6248_1562# vdd.t528 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X299 swmatrix_Tgate_2.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t295 vss.t294 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X300 BUS[6].t9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t96 vdd.t236 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X301 pin.t224 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 BUS[1].t18 vdd.t518 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X302 BUS[4].t9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t193 vdd.t439 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X303 swmatrix_Tgate_6.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t382 vdd.t381 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X304 a_54841_1539# ShiftReg_row_10_2$1_0.Q[9] vss.t6 vss.t5 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X305 a_9696_2122# a_8712_1562# a_9548_2122# vdd.t419 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X306 pin.t197 swmatrix_Tgate_9.gated_control BUS[1].t14 vss.t339 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X307 a_41100_2122# a_40380_1580# a_40896_2122# vdd.t23 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X308 vdd.t386 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] vdd.t385 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X309 BUS[1].t19 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 pin.t225 vdd.t519 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X310 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[7] vdd.t390 vdd.t389 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X311 a_19712_2122# a_19196_1580# a_19564_1577# vss.t75 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X312 pin.t55 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[8].t9 vdd.t116 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X313 a_3800_2002# a_3456_2122# vss.t203 vss.t202 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X314 vdd.t192 a_10040_2002# a_9900_2122# vdd.t191 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X315 a_59100_1580# a_58632_1562# vss.t313 vss.t312 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X316 vdd.t255 phi_2.t9 a_8712_1562# vdd.t254 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X317 pin.t213 swmatrix_Tgate_0.gated_control BUS[7].t18 vss.t388 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X318 a_47136_2122# a_46152_1562# a_46988_2122# vdd.t437 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X319 vss.t230 a_32536_2002# a_32436_1577# vss.t229 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X320 BUS[10].t21 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 pin.t166 vdd.t367 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X321 a_1236_1577# a_8_1562# a_992_2122# vss.t2 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X322 BUS[7].t10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 pin.t92 vdd.t232 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X323 BUS[4].t8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 pin.t128 vdd.t308 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X324 a_31676_1580# a_31208_1562# vss.t99 vss.t98 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X325 vdd.t239 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t238 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X326 vss.t49 phi_1.t10 a_43688_1562# vss.t48 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X327 a_38776_2002# a_38432_2122# vss.t139 vss.t138 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X328 a_59960_2002# a_59616_2122# vdd.t217 vdd.t216 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X329 a_50396_1580# a_49928_1562# vdd.t144 vdd.t143 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X330 pin.t111 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 BUS[10].t10 vdd.t276 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X331 a_53720_2002# a_53376_2122# vdd.t384 vdd.t383 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X332 a_13676_2122# a_12956_1580# a_13472_2122# vdd.t515 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X333 pin.t97 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[6].t8 vdd.t237 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X334 BUS[3].t4 swmatrix_Tgate_4.gated_control pin.t173 vss.t261 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X335 pin.t43 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[2].t5 vdd.t105 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X336 pin.t129 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 BUS[4].t7 vdd.t309 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X337 swmatrix_Tgate_8.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t65 vdd.t64 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X338 pin.t121 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[9].t3 vdd.t295 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X339 vss.t192 phi_2.t10 a_14952_1562# vss.t191 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X340 vdd.t393 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t392 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X341 vdd.t453 a_1336_2002# a_1196_2122# vdd.t452 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X342 pin.t172 swmatrix_Tgate_4.gated_control BUS[3].t3 vss.t260 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X343 BUS[2].t4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 pin.t8 vdd.t24 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X344 vss.t225 a_41240_2002# a_41140_1577# vss.t224 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X345 a_15420_1580# a_14952_1562# vdd.t330 vdd.t329 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X346 pin.t226 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 BUS[1].t20 vdd.t520 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X347 a_40380_1580# a_39912_1562# vss.t293 vss.t292 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X348 pin.t203 swmatrix_Tgate_7.gated_control BUS[4].t20 vss.t367 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X349 BUS[7].t9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 pin.t222 vdd.t513 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X350 vss.t208 phi_2.t11 a_52392_1562# vss.t207 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X351 a_19712_2122# a_18728_1562# a_19564_2122# vdd.t158 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X352 BUS[3].t12 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 pin.t101 vdd.t247 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X353 a_22380_2122# a_21660_1580# a_22176_2122# vdd.t180 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X354 BUS[10].t11 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 pin.t112 vdd.t277 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X355 a_52860_1580# a_52392_1562# vdd.t279 vdd.t278 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X356 a_38676_1577# a_37448_1562# a_38432_2122# vss.t226 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X357 vss.t53 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t52 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X358 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t10 a_61081_1539# vss.t355 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X359 pin.t223 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[7].t8 vdd.t514 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X360 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t11 a_54841_1539# vss.t344 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X361 a_19564_1577# ShiftReg_row_10_2$1_0.Q[3] vss.t402 vss.t401 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X362 pin.t37 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 BUS[5].t8 vdd.t80 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X363 vss.t338 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t337 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X364 vdd.t67 phi_1.t11 a_24968_1562# vdd.t66 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X365 a_32536_2002# a_32192_2122# vdd.t376 vdd.t375 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X366 pin.t102 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[3].t11 vdd.t248 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X367 vdd.t69 phi_1.t12 a_18728_1562# vdd.t68 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X368 vdd.t458 enable.t12 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t457 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X369 vdd.t413 a_3800_2002# a_3660_2122# vdd.t412 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X370 pin.t178 swmatrix_Tgate_6.gated_control BUS[6].t20 vss.t281 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X371 vss.t239 phi_1.t13 a_6248_1562# vss.t238 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X372 BUS[1].t13 swmatrix_Tgate_9.gated_control pin.t196 vss.t336 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X373 a_57004_1577# ShiftReg_row_10_2$1_0.Q[9] vss.t4 vss.t3 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X374 BUS[5].t7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 pin.t32 vdd.t79 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X375 a_40896_2122# a_40380_1580# a_40748_1577# vss.t14 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X376 a_6716_1580# a_6248_1562# vdd.t369 vdd.t368 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X377 a_51256_2002# a_50912_2122# vss.t164 vss.t163 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X378 a_7084_2122# ShiftReg_row_10_2$1_0.Q[1] vdd.t447 vdd.t446 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X379 vdd.t372 a_38776_2002# a_38636_2122# vdd.t371 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X380 BUS[6].t7 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 pin.t98 vdd.t244 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X381 a_47380_1577# a_46152_1562# a_47136_2122# vss.t316 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X382 a_16280_2002# a_15936_2122# vss.t83 vss.t82 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X383 BUS[10].t2 swmatrix_Tgate_2.gated_control pin.t49 vss.t69 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X384 a_476_1580# a_8_1562# vss.t1 vss.t0 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X385 BUS[8].t4 swmatrix_Tgate_3.gated_control pin.t12 vss.t19 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X386 vss.t137 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t136 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X387 swmatrix_Tgate_9.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t146 vss.t145 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X388 vdd.t290 phi_2.t12 a_27432_1562# vdd.t289 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X389 pin.t184 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[8].t19 vdd.t407 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X390 vdd.t177 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] vdd.t176 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X391 pin.t48 swmatrix_Tgate_2.gated_control BUS[10].t1 vss.t68 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X392 a_53720_2002# a_53376_2122# vss.t268 vss.t267 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X393 vss.t210 phi_2.t13 a_8712_1562# vss.t209 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X394 a_44524_2122# ShiftReg_row_10_2$1_0.Q[7] vdd.t388 vdd.t387 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X395 vss.t387 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t386 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X396 a_59616_2122# a_59100_1580# a_59468_1577# vss.t343 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X397 vdd.t460 enable.t13 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t459 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X398 BUS[5].t6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 pin.t30 vdd.t78 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X399 vdd.t307 a_47480_2002# a_47340_2122# vdd.t306 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X400 BUS[2].t3 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 pin.t9 vdd.t25 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X401 a_51116_2122# a_50396_1580# a_50912_2122# vdd.t141 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X402 BUS[2].t20 swmatrix_Tgate_8.gated_control pin.t68 vss.t122 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X403 a_32044_1577# ShiftReg_row_10_2$1_0.Q[5] vss.t130 vss.t129 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X404 vss.t170 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] vss.t169 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X405 a_36121_1539# ShiftReg_row_10_2$1_0.Q[6] vss.t216 vss.t215 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X406 pin.t33 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[5].t5 vdd.t77 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X407 vdd.t503 a_20056_2002# a_19916_2122# vdd.t502 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X408 a_3456_2122# a_2940_1580# a_3308_1577# vss.t176 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X409 vdd.t488 a_13816_2002# a_13676_2122# vdd.t487 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X410 a_46988_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t182 vdd.t181 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X411 a_22420_1577# a_21192_1562# a_22176_2122# vss.t193 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X412 a_40896_2122# a_39912_1562# a_40748_2122# vdd.t404 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X413 pin.t66 swmatrix_Tgate_8.gated_control BUS[2].t19 vss.t121 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X414 pin.t70 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[4].t6 vdd.t183 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X415 pin.t227 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[1].t21 vdd.t521 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X416 vdd.t128 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t127 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X417 BUS[8].t20 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 pin.t185 vdd.t408 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X418 BUS[6].t6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 pin.t99 vdd.t245 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X419 a_38432_2122# a_37916_1580# a_38284_1577# vss.t142 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X420 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[9] vdd.t12 vdd.t11 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X421 pin.t83 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[10].t8 vdd.t223 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X422 pin.t186 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[8].t21 vdd.t409 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X423 vdd.t162 a_22520_2002# a_22380_2122# vdd.t161 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X424 pin.t100 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[6].t5 vdd.t246 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X425 vss.t241 phi_1.t14 a_24968_1562# vss.t240 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X426 vss.t243 phi_1.t15 a_18728_1562# vss.t242 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X427 a_59616_2122# a_58632_1562# a_59468_2122# vdd.t432 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X428 a_35000_2002# a_34656_2122# vdd.t479 vdd.t478 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X429 pin.t144 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 BUS[7].t7 vdd.t324 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X430 vss.t51 a_51256_2002# a_51156_1577# vss.t50 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X431 a_25436_1580# a_24968_1562# vdd.t417 vdd.t416 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X432 BUS[2].t2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 pin.t75 vdd.t193 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X433 a_50396_1580# a_49928_1562# vss.t103 vss.t102 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X434 BUS[4].t5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 pin.t132 vdd.t312 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X435 pin.t228 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[1].t22 vdd.t522 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X436 a_22028_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t171 vdd.t170 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X437 vss.t280 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t279 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X438 BUS[9].t11 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 pin.t160 vdd.t357 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X439 a_59468_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t394 vss.t393 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X440 a_32396_2122# a_31676_1580# a_32192_2122# vdd.t338 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X441 swmatrix_Tgate_7.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t77 vss.t76 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X442 swmatrix_Tgate_5.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t126 vdd.t125 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X443 pin.t145 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[7].t6 vdd.t325 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X444 BUS[4].t19 swmatrix_Tgate_7.gated_control pin.t202 vss.t366 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X445 a_3456_2122# a_2472_1562# a_3308_2122# vdd.t97 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X446 a_9548_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t52 vdd.t51 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X447 vss.t94 a_16280_2002# a_16180_1577# vss.t93 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X448 pin.t76 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[2].t1 vdd.t194 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X449 swmatrix_Tgate_4.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t79 vss.t78 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X450 BUS[1].t9 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 pin.t118 vdd.t286 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X451 a_15420_1580# a_14952_1562# vss.t222 vss.t221 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X452 vss.t245 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] vss.t244 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X453 a_17401_1539# ShiftReg_row_10_2$1_0.Q[3] vss.t400 vss.t399 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X454 pin.t72 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 BUS[8].t10 vdd.t185 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X455 pin.t161 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 BUS[9].t12 vdd.t358 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X456 pin.t181 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 BUS[6].t4 vdd.t394 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X457 BUS[3].t2 swmatrix_Tgate_4.gated_control pin.t171 vss.t259 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X458 vss.t212 phi_2.t14 a_27432_1562# vss.t211 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X459 a_844_1577# D_in.t1 vss.t405 vss.t404 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X460 a_3308_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t332 vss.t331 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X461 a_34140_1580# a_33672_1562# vdd.t190 vdd.t189 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X462 pin.t103 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 BUS[3].t10 vdd.t249 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X463 vss.t40 a_53720_2002# a_53620_1577# vss.t39 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X464 a_27900_1580# a_27432_1562# vdd.t132 vdd.t131 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X465 pin.t84 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 BUS[10].t9 vdd.t224 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X466 vdd.t27 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t26 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X467 a_52860_1580# a_52392_1562# vss.t205 vss.t204 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X468 pin.t58 swmatrix_Tgate_5.gated_control BUS[5].t19 vss.t113 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X469 a_38432_2122# a_37448_1562# a_38284_2122# vdd.t335 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X470 BUS[8].t11 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 pin.t73 vdd.t186 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X471 a_13816_2002# a_13472_2122# vdd.t29 vdd.t28 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X472 a_50912_2122# a_50396_1580# a_50764_1577# vss.t100 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X473 a_34860_2122# a_34140_1580# a_34656_2122# vdd.t429 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X474 a_57396_1577# a_56168_1562# a_57152_2122# vss.t351 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X475 BUS[7].t5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 pin.t149 vdd.t342 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X476 BUS[7].t17 swmatrix_Tgate_0.gated_control pin.t218 vss.t385 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X477 pin.t127 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[10].t12 vdd.t305 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X478 a_22176_2122# a_21660_1580# a_22028_1577# vss.t153 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X479 a_38284_1577# ShiftReg_row_10_2$1_0.Q[6] vss.t214 vss.t213 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X480 vss.t182 a_7576_2002# a_7476_1577# vss.t181 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X481 a_15936_2122# a_15420_1580# a_15788_1577# vss.t96 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X482 vdd.t301 phi_1.t16 a_37448_1562# vdd.t300 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X483 a_51256_2002# a_50912_2122# vdd.t197 vdd.t196 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X484 pin.t36 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 BUS[5].t4 vdd.t76 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X485 vdd.t467 enable.t14 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t466 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X486 pin.t155 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 BUS[9].t9 vdd.t352 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X487 vdd.t90 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t89 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X488 pin.t150 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 BUS[7].t4 vdd.t347 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X489 a_16280_2002# a_15936_2122# vdd.t122 vdd.t121 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X490 vdd.t485 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t484 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X491 pin.t11 swmatrix_Tgate_3.gated_control BUS[8].t3 vss.t18 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X492 BUS[9].t10 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 pin.t156 vdd.t353 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X493 vdd.t211 a_57496_2002# a_57356_2122# vdd.t210 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X494 BUS[3].t9 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 pin.t93 vdd.t233 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X495 a_59860_1577# a_58632_1562# a_59616_2122# vss.t311 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X496 a_35000_2002# a_34656_2122# vss.t357 vss.t356 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X497 BUS[10].t13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 pin.t138 vdd.t318 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X498 vss.t285 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] vss.t284 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X499 BUS[10].t0 swmatrix_Tgate_2.gated_control pin.t47 vss.t67 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X500 vss.t64 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t63 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X501 vdd.t33 phi_2.t15 a_46152_1562# vdd.t32 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X502 pin.t41 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[5].t3 vdd.t75 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X503 a_32436_1577# a_31208_1562# a_32192_2122# vss.t97 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X504 pin.t94 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 BUS[3].t8 vdd.t234 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X505 pin.t139 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[10].t14 vdd.t319 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X506 vdd.t164 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t163 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X507 a_3700_1577# a_2472_1562# a_3456_2122# vss.t60 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X508 a_13324_1577# ShiftReg_row_10_2$1_0.Q[2] vss.t32 vss.t31 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X509 pin.t65 swmatrix_Tgate_8.gated_control BUS[2].t18 vss.t120 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X510 a_57004_2122# ShiftReg_row_10_2$1_0.Q[9] vdd.t10 vdd.t9 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X511 a_50912_2122# a_49928_1562# a_50764_2122# vdd.t142 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X512 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t15 a_17401_1539# vss.t347 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X513 vdd.t469 enable.t16 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t468 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X514 BUS[5].t2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 pin.t29 vdd.t74 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X515 vdd.t524 a_59960_2002# a_59820_2122# vdd.t523 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X516 a_28268_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t209 vdd.t208 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X517 a_22176_2122# a_21192_1562# a_22028_2122# vdd.t258 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X518 a_15936_2122# a_14952_1562# a_15788_2122# vdd.t328 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X519 a_50764_1577# ShiftReg_row_10_2$1_0.Q[8] vss.t320 vss.t319 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X520 BUS[2].t17 swmatrix_Tgate_8.gated_control pin.t64 vss.t119 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X521 BUS[4].t4 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 pin.t133 vdd.t313 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X522 vdd.t337 a_32536_2002# a_32396_2122# vdd.t336 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X523 a_13816_2002# a_13472_2122# vss.t26 vss.t25 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X524 pin.t164 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[9].t13 vdd.t365 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X525 BUS[6].t19 swmatrix_Tgate_6.gated_control pin.t177 vss.t278 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X526 a_41140_1577# a_39912_1562# a_40896_2122# vss.t291 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X527 a_15788_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t349 vss.t348 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X528 a_10040_2002# a_9696_2122# vss.t148 vss.t147 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X529 pin.t182 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[6].t3 vdd.t395 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X530 BUS[1].t10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 pin.t119 vdd.t287 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X531 vdd.t205 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] vdd.t204 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X532 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[6] vdd.t292 vdd.t291 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X533 pin.t167 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[4].t3 vdd.t373 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X534 vdd.t35 phi_2.t16 a_21192_1562# vdd.t34 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X535 pin.t10 swmatrix_Tgate_3.gated_control BUS[8].t2 vss.t17 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X536 vss.t201 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] vss.t200 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X537 BUS[3].t7 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 pin.t95 vdd.t235 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X538 pin.t120 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 BUS[1].t11 vdd.t288 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X539 a_57152_2122# a_56636_1580# a_57004_1577# vss.t350 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X540 vss.t382 a_26296_2002# a_26196_1577# vss.t381 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X541 vdd.t332 a_41240_2002# a_41100_2122# vdd.t331 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X542 a_25436_1580# a_24968_1562# vss.t299 vss.t298 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X543 pin.t28 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[5].t1 vdd.t73 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X544 vss.t218 phi_1.t17 a_37448_1562# vss.t217 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X545 BUS[9].t17 swmatrix_Tgate_1.gated_control pin.t207 vss.t374 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X546 pin.t71 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[3].t6 vdd.t184 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X547 a_13716_1577# a_12488_1562# a_13472_2122# vss.t41 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X548 a_44156_1580# a_43688_1562# vdd.t148 vdd.t147 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X549 a_37916_1580# a_37448_1562# vdd.t334 vdd.t333 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X550 pin.t168 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 BUS[4].t2 vdd.t374 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X551 pin.t201 swmatrix_Tgate_7.gated_control BUS[4].t18 vss.t365 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X552 pin.t82 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[2].t0 vdd.t220 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X553 a_40748_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t179 vdd.t178 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X554 BUS[6].t2 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 pin.t183 vdd.t396 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X555 pin.t170 swmatrix_Tgate_4.gated_control BUS[3].t1 vss.t258 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X556 a_44876_2122# a_44156_1580# a_44672_2122# vdd.t63 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X557 vss.t57 a_35000_2002# a_34900_1577# vss.t56 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X558 BUS[4].t1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 pin.t141 vdd.t321 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X559 pin.t50 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[1].t3 vdd.t108 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X560 vss.t59 a_28760_2002# a_28660_1577# vss.t58 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X561 swmatrix_Tgate_6.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t266 vss.t265 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X562 vss.t16 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t15 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X563 swmatrix_Tgate_0.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t506 vdd.t505 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X564 a_34140_1580# a_33672_1562# vss.t157 vss.t156 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X565 a_29881_1539# ShiftReg_row_10_2$1_0.Q[5] vss.t128 vss.t127 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X566 vss.t28 phi_2.t17 a_46152_1562# vss.t27 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X567 pin.t74 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[8].t12 vdd.t187 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X568 BUS[5].t18 swmatrix_Tgate_5.gated_control pin.t62 vss.t112 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X569 a_992_2122# a_476_1580# a_844_1577# vss.t346 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X570 pin.t116 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[6].t1 vdd.t284 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X571 BUS[1].t4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 pin.t51 vdd.t109 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X572 a_46620_1580# a_46152_1562# vdd.t436 vdd.t435 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X573 a_7576_2002# a_7232_2122# vss.t184 vss.t183 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X574 a_16140_2122# a_15420_1580# a_15936_2122# vdd.t137 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X575 vdd.t364 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] vdd.t363 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X576 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I ShiftReg_row_10_2$1_0.Q[3] vdd.t510 vdd.t509 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X577 vss.t24 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t23 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X578 pin.t151 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 BUS[7].t3 vdd.t348 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X579 vdd.t107 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t106 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X580 a_57152_2122# a_56168_1562# a_57004_2122# vdd.t473 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X581 a_26296_2002# a_25952_2122# vdd.t424 vdd.t423 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X582 a_53580_2122# a_52860_1580# a_53376_2122# vdd.t403 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X583 BUS[10].t15 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 pin.t146 vdd.t326 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X584 vss.t364 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss.t363 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X585 vss.t162 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t161 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X586 BUS[7].t2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 pin.t122 vdd.t296 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X587 a_34656_2122# a_34140_1580# a_34508_1577# vss.t310 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X588 vdd.t303 phi_1.t18 a_56168_1562# vdd.t302 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X589 a_53228_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss.t166 vss.t165 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X590 BUS[9].t16 swmatrix_Tgate_1.gated_control pin.t206 vss.t373 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X591 a_3308_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t451 vdd.t450 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X592 pin.t134 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 BUS[9].t6 vdd.t314 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X593 swmatrix_Tgate_8.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss.t47 vss.t46 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X594 pin.t107 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[4].t0 vdd.t264 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X595 vss.t36 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] vss.t35 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X596 a_28760_2002# a_28416_2122# vdd.t362 vdd.t361 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X597 a_7436_2122# a_6716_1580# a_7232_2122# vdd.t136 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X598 a_11161_1539# ShiftReg_row_10_2$1_0.Q[2] vss.t30 vss.t29 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X599 vss.t81 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] vss.t80 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X600 vdd.t153 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t152 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X601 pin.t169 swmatrix_Tgate_4.gated_control BUS[3].t0 vss.t257 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X602 BUS[6].t0 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 pin.t117 vdd.t285 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X603 vss.t178 a_59616_2122# d_out.t0 vss.t177 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X604 a_47480_2002# a_47136_2122# vss.t168 vss.t167 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X605 a_992_2122# a_8_1562# a_844_2122# vdd.t6 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X606 BUS[7].t1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 pin.t123 vdd.t297 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X607 vdd.t37 phi_2.t18 a_58632_1562# vdd.t36 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X608 BUS[5].t17 swmatrix_Tgate_5.gated_control pin.t63 vss.t111 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X609 a_51156_1577# a_49928_1562# a_50912_2122# vss.t101 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X610 vdd.t398 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] vdd.t397 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X611 a_13472_2122# a_12956_1580# a_13324_1577# vss.t403 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X612 vdd.t101 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd.t100 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X613 pin.t135 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 BUS[9].t7 vdd.t315 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X614 BUS[6].t18 swmatrix_Tgate_6.gated_control pin.t176 vss.t277 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X615 pin.t219 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[7].t0 vdd.t504 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X616 BUS[4].t17 swmatrix_Tgate_7.gated_control pin.t200 vss.t362 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X617 vdd.t257 phi_1.t19 a_31208_1562# vdd.t256 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X618 a_9900_2122# a_9180_1580# a_9696_2122# vdd.t212 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X619 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t17 a_36121_1539# vss.t360 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X620 pin.t39 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 BUS[5].t0 vdd.t72 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X621 vdd.t483 enable.t18 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd.t482 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X622 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable.t19 a_29881_1539# vss.t361 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X623 vdd.t243 phi_2.t19 a_2472_1562# vdd.t242 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X624 vdd.t490 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vdd.t489 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X625 a_10040_2002# a_9696_2122# vdd.t175 vdd.t174 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X626 a_34656_2122# a_33672_1562# a_34508_2122# vdd.t188 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X627 BUS[9].t2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 pin.t108 vdd.t273 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X628 pin.t175 swmatrix_Tgate_6.gated_control BUS[6].t17 vss.t276 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X629 BUS[1].t12 swmatrix_Tgate_9.gated_control pin.t195 vss.t335 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
R0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.7994
R1 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R3 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R4 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R5 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R11 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R13 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R17 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R18 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R19 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R20 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R21 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R22 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R23 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R24 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R25 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R26 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R27 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R28 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R29 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R30 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R31 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R32 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R33 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R34 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R35 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R36 pin.n100 pin.t84 11.5207
R37 pin.n108 pin.t44 11.3417
R38 pin.n111 pin.t49 11.3417
R39 pin.n121 pin.t211 11.3417
R40 pin.n124 pin.t206 11.3417
R41 pin.n134 pin.t11 11.3417
R42 pin.n137 pin.t13 11.3417
R43 pin.n147 pin.t213 11.3417
R44 pin.n150 pin.t217 11.3417
R45 pin.n160 pin.t178 11.3417
R46 pin.n163 pin.t176 11.3417
R47 pin.n173 pin.t61 11.3417
R48 pin.n176 pin.t63 11.3417
R49 pin.n186 pin.t204 11.3417
R50 pin.n189 pin.t202 11.3417
R51 pin.n199 pin.t170 11.3417
R52 pin.n202 pin.t173 11.3417
R53 pin.n212 pin.t69 11.3417
R54 pin.n215 pin.t68 11.3417
R55 pin.n225 pin.t194 11.3417
R56 pin.n228 pin.t198 11.3417
R57 pin.n112 pin.t161 11.2907
R58 pin.n125 pin.t54 11.2907
R59 pin.n138 pin.t126 11.2907
R60 pin.n151 pin.t212 11.2907
R61 pin.n164 pin.t36 11.2907
R62 pin.n177 pin.t167 11.2907
R63 pin.n190 pin.t102 11.2907
R64 pin.n203 pin.t56 11.2907
R65 pin.n216 pin.t18 11.2907
R66 pin.n109 pin.n91 10.7117
R67 pin.n110 pin.n90 10.7117
R68 pin.n122 pin.n81 10.7117
R69 pin.n123 pin.n80 10.7117
R70 pin.n135 pin.n71 10.7117
R71 pin.n136 pin.n70 10.7117
R72 pin.n148 pin.n61 10.7117
R73 pin.n149 pin.n60 10.7117
R74 pin.n161 pin.n51 10.7117
R75 pin.n162 pin.n50 10.7117
R76 pin.n174 pin.n41 10.7117
R77 pin.n175 pin.n40 10.7117
R78 pin.n187 pin.n31 10.7117
R79 pin.n188 pin.n30 10.7117
R80 pin.n200 pin.n21 10.7117
R81 pin.n201 pin.n20 10.7117
R82 pin.n213 pin.n11 10.7117
R83 pin.n214 pin.n10 10.7117
R84 pin.n226 pin.n1 10.7117
R85 pin.n227 pin.n0 10.7117
R86 pin.n100 pin.n99 10.5557
R87 pin.n101 pin.n98 10.5557
R88 pin.n102 pin.n97 10.5557
R89 pin.n103 pin.n96 10.5557
R90 pin.n104 pin.n95 10.5557
R91 pin.n105 pin.n94 10.5557
R92 pin.n106 pin.n93 10.5557
R93 pin.n107 pin.n92 10.5557
R94 pin.n113 pin.n89 10.5557
R95 pin.n114 pin.n88 10.5557
R96 pin.n115 pin.n87 10.5557
R97 pin.n116 pin.n86 10.5557
R98 pin.n117 pin.n85 10.5557
R99 pin.n118 pin.n84 10.5557
R100 pin.n119 pin.n83 10.5557
R101 pin.n120 pin.n82 10.5557
R102 pin.n126 pin.n79 10.5557
R103 pin.n127 pin.n78 10.5557
R104 pin.n128 pin.n77 10.5557
R105 pin.n129 pin.n76 10.5557
R106 pin.n130 pin.n75 10.5557
R107 pin.n131 pin.n74 10.5557
R108 pin.n132 pin.n73 10.5557
R109 pin.n133 pin.n72 10.5557
R110 pin.n139 pin.n69 10.5557
R111 pin.n140 pin.n68 10.5557
R112 pin.n141 pin.n67 10.5557
R113 pin.n142 pin.n66 10.5557
R114 pin.n143 pin.n65 10.5557
R115 pin.n144 pin.n64 10.5557
R116 pin.n145 pin.n63 10.5557
R117 pin.n146 pin.n62 10.5557
R118 pin.n152 pin.n59 10.5557
R119 pin.n153 pin.n58 10.5557
R120 pin.n154 pin.n57 10.5557
R121 pin.n155 pin.n56 10.5557
R122 pin.n156 pin.n55 10.5557
R123 pin.n157 pin.n54 10.5557
R124 pin.n158 pin.n53 10.5557
R125 pin.n159 pin.n52 10.5557
R126 pin.n165 pin.n49 10.5557
R127 pin.n166 pin.n48 10.5557
R128 pin.n167 pin.n47 10.5557
R129 pin.n168 pin.n46 10.5557
R130 pin.n169 pin.n45 10.5557
R131 pin.n170 pin.n44 10.5557
R132 pin.n171 pin.n43 10.5557
R133 pin.n172 pin.n42 10.5557
R134 pin.n178 pin.n39 10.5557
R135 pin.n179 pin.n38 10.5557
R136 pin.n180 pin.n37 10.5557
R137 pin.n181 pin.n36 10.5557
R138 pin.n182 pin.n35 10.5557
R139 pin.n183 pin.n34 10.5557
R140 pin.n184 pin.n33 10.5557
R141 pin.n185 pin.n32 10.5557
R142 pin.n191 pin.n29 10.5557
R143 pin.n192 pin.n28 10.5557
R144 pin.n193 pin.n27 10.5557
R145 pin.n194 pin.n26 10.5557
R146 pin.n195 pin.n25 10.5557
R147 pin.n196 pin.n24 10.5557
R148 pin.n197 pin.n23 10.5557
R149 pin.n198 pin.n22 10.5557
R150 pin.n204 pin.n19 10.5557
R151 pin.n205 pin.n18 10.5557
R152 pin.n206 pin.n17 10.5557
R153 pin.n207 pin.n16 10.5557
R154 pin.n208 pin.n15 10.5557
R155 pin.n209 pin.n14 10.5557
R156 pin.n210 pin.n13 10.5557
R157 pin.n211 pin.n12 10.5557
R158 pin.n217 pin.n9 10.5557
R159 pin.n218 pin.n8 10.5557
R160 pin.n219 pin.n7 10.5557
R161 pin.n220 pin.n6 10.5557
R162 pin.n221 pin.n5 10.5557
R163 pin.n222 pin.n4 10.5557
R164 pin.n223 pin.n3 10.5557
R165 pin.n224 pin.n2 10.5557
R166 pin.n216 pin 0.731668
R167 pin.n112 pin 0.67123
R168 pin.n125 pin 0.67123
R169 pin.n138 pin 0.67123
R170 pin.n151 pin 0.67123
R171 pin.n164 pin 0.67123
R172 pin.n177 pin 0.67123
R173 pin.n190 pin 0.67123
R174 pin.n203 pin 0.67123
R175 pin pin.n111 0.564807
R176 pin pin.n124 0.564807
R177 pin pin.n137 0.564807
R178 pin pin.n150 0.564807
R179 pin pin.n163 0.564807
R180 pin pin.n176 0.564807
R181 pin pin.n189 0.564807
R182 pin pin.n202 0.564807
R183 pin pin.n215 0.564807
R184 pin pin.n228 0.564807
R185 pin.n108 pin.n107 0.496485
R186 pin.n121 pin.n120 0.496485
R187 pin.n134 pin.n133 0.496485
R188 pin.n147 pin.n146 0.496485
R189 pin.n160 pin.n159 0.496485
R190 pin.n173 pin.n172 0.496485
R191 pin.n186 pin.n185 0.496485
R192 pin.n199 pin.n198 0.496485
R193 pin.n212 pin.n211 0.496485
R194 pin.n225 pin.n224 0.496485
R195 pin.n99 pin.t112 0.4555
R196 pin.n99 pin.t158 0.4555
R197 pin.n98 pin.t162 0.4555
R198 pin.n98 pin.t139 0.4555
R199 pin.n97 pin.t157 0.4555
R200 pin.n97 pin.t189 0.4555
R201 pin.n96 pin.t138 0.4555
R202 pin.n96 pin.t111 0.4555
R203 pin.n95 pin.t80 0.4555
R204 pin.n95 pin.t83 0.4555
R205 pin.n94 pin.t166 0.4555
R206 pin.n94 pin.t147 0.4555
R207 pin.n93 pin.t146 0.4555
R208 pin.n93 pin.t127 0.4555
R209 pin.n92 pin.t163 0.4555
R210 pin.n92 pin.t81 0.4555
R211 pin.n89 pin.t78 0.4555
R212 pin.n89 pin.t124 0.4555
R213 pin.n88 pin.t160 0.4555
R214 pin.n88 pin.t121 0.4555
R215 pin.n87 pin.t148 0.4555
R216 pin.n87 pin.t134 0.4555
R217 pin.n86 pin.t156 0.4555
R218 pin.n86 pin.t187 0.4555
R219 pin.n85 pin.t221 0.4555
R220 pin.n85 pin.t155 0.4555
R221 pin.n84 pin.t79 0.4555
R222 pin.n84 pin.t125 0.4555
R223 pin.n83 pin.t108 0.4555
R224 pin.n83 pin.t164 0.4555
R225 pin.n82 pin.t188 0.4555
R226 pin.n82 pin.t135 0.4555
R227 pin.n79 pin.t6 0.4555
R228 pin.n79 pin.t184 0.4555
R229 pin.n78 pin.t106 0.4555
R230 pin.n78 pin.t229 0.4555
R231 pin.n77 pin.t113 0.4555
R232 pin.n77 pin.t186 0.4555
R233 pin.n76 pin.t115 0.4555
R234 pin.n76 pin.t7 0.4555
R235 pin.n75 pin.t185 0.4555
R236 pin.n75 pin.t55 0.4555
R237 pin.n74 pin.t105 0.4555
R238 pin.n74 pin.t74 0.4555
R239 pin.n73 pin.t73 0.4555
R240 pin.n73 pin.t104 0.4555
R241 pin.n72 pin.t114 0.4555
R242 pin.n72 pin.t72 0.4555
R243 pin.n69 pin.t165 0.4555
R244 pin.n69 pin.t144 0.4555
R245 pin.n68 pin.t92 0.4555
R246 pin.n68 pin.t137 0.4555
R247 pin.n67 pin.t122 0.4555
R248 pin.n67 pin.t150 0.4555
R249 pin.n66 pin.t136 0.4555
R250 pin.n66 pin.t151 0.4555
R251 pin.n65 pin.t149 0.4555
R252 pin.n65 pin.t223 0.4555
R253 pin.n64 pin.t110 0.4555
R254 pin.n64 pin.t219 0.4555
R255 pin.n63 pin.t222 0.4555
R256 pin.n63 pin.t109 0.4555
R257 pin.n62 pin.t123 0.4555
R258 pin.n62 pin.t145 0.4555
R259 pin.n59 pin.t98 0.4555
R260 pin.n59 pin.t100 0.4555
R261 pin.n58 pin.t22 0.4555
R262 pin.n58 pin.t182 0.4555
R263 pin.n57 pin.t99 0.4555
R264 pin.n57 pin.t154 0.4555
R265 pin.n56 pin.t152 0.4555
R266 pin.n56 pin.t116 0.4555
R267 pin.n55 pin.t96 0.4555
R268 pin.n55 pin.t24 0.4555
R269 pin.n54 pin.t183 0.4555
R270 pin.n54 pin.t181 0.4555
R271 pin.n53 pin.t23 0.4555
R272 pin.n53 pin.t153 0.4555
R273 pin.n52 pin.t117 0.4555
R274 pin.n52 pin.t97 0.4555
R275 pin.n49 pin.t32 0.4555
R276 pin.n49 pin.t27 0.4555
R277 pin.n48 pin.t25 0.4555
R278 pin.n48 pin.t37 0.4555
R279 pin.n47 pin.t31 0.4555
R280 pin.n47 pin.t39 0.4555
R281 pin.n46 pin.t29 0.4555
R282 pin.n46 pin.t33 0.4555
R283 pin.n45 pin.t40 0.4555
R284 pin.n45 pin.t41 0.4555
R285 pin.n44 pin.t30 0.4555
R286 pin.n44 pin.t26 0.4555
R287 pin.n43 pin.t34 0.4555
R288 pin.n43 pin.t28 0.4555
R289 pin.n42 pin.t38 0.4555
R290 pin.n42 pin.t35 0.4555
R291 pin.n39 pin.t140 0.4555
R292 pin.n39 pin.t130 0.4555
R293 pin.n38 pin.t133 0.4555
R294 pin.n38 pin.t70 0.4555
R295 pin.n37 pin.t193 0.4555
R296 pin.n37 pin.t159 0.4555
R297 pin.n36 pin.t141 0.4555
R298 pin.n36 pin.t192 0.4555
R299 pin.n35 pin.t131 0.4555
R300 pin.n35 pin.t168 0.4555
R301 pin.n34 pin.t132 0.4555
R302 pin.n34 pin.t129 0.4555
R303 pin.n33 pin.t143 0.4555
R304 pin.n33 pin.t107 0.4555
R305 pin.n32 pin.t128 0.4555
R306 pin.n32 pin.t142 0.4555
R307 pin.n29 pin.t19 0.4555
R308 pin.n29 pin.t103 0.4555
R309 pin.n28 pin.t101 0.4555
R310 pin.n28 pin.t91 0.4555
R311 pin.n27 pin.t21 0.4555
R312 pin.n27 pin.t94 0.4555
R313 pin.n26 pin.t90 0.4555
R314 pin.n26 pin.t20 0.4555
R315 pin.n25 pin.t93 0.4555
R316 pin.n25 pin.t71 0.4555
R317 pin.n24 pin.t191 0.4555
R318 pin.n24 pin.t52 0.4555
R319 pin.n23 pin.t95 0.4555
R320 pin.n23 pin.t190 0.4555
R321 pin.n22 pin.t89 0.4555
R322 pin.n22 pin.t53 0.4555
R323 pin.n19 pin.t3 0.4555
R324 pin.n19 pin.t77 0.4555
R325 pin.n18 pin.t9 0.4555
R326 pin.n18 pin.t42 0.4555
R327 pin.n17 pin.t220 0.4555
R328 pin.n17 pin.t82 0.4555
R329 pin.n16 pin.t57 0.4555
R330 pin.n16 pin.t4 0.4555
R331 pin.n15 pin.t1 0.4555
R332 pin.n15 pin.t76 0.4555
R333 pin.n14 pin.t8 0.4555
R334 pin.n14 pin.t0 0.4555
R335 pin.n13 pin.t75 0.4555
R336 pin.n13 pin.t43 0.4555
R337 pin.n12 pin.t5 0.4555
R338 pin.n12 pin.t2 0.4555
R339 pin.n9 pin.t88 0.4555
R340 pin.n9 pin.t120 0.4555
R341 pin.n8 pin.t17 0.4555
R342 pin.n8 pin.t16 0.4555
R343 pin.n7 pin.t119 0.4555
R344 pin.n7 pin.t227 0.4555
R345 pin.n6 pin.t225 0.4555
R346 pin.n6 pin.t86 0.4555
R347 pin.n5 pin.t51 0.4555
R348 pin.n5 pin.t224 0.4555
R349 pin.n4 pin.t85 0.4555
R350 pin.n4 pin.t50 0.4555
R351 pin.n3 pin.t118 0.4555
R352 pin.n3 pin.t226 0.4555
R353 pin.n2 pin.t87 0.4555
R354 pin.n2 pin.t228 0.4555
R355 pin.n91 pin.t47 0.41
R356 pin.n91 pin.t48 0.41
R357 pin.n90 pin.t45 0.41
R358 pin.n90 pin.t46 0.41
R359 pin.n81 pin.t207 0.41
R360 pin.n81 pin.t210 0.41
R361 pin.n80 pin.t208 0.41
R362 pin.n80 pin.t209 0.41
R363 pin.n71 pin.t12 0.41
R364 pin.n71 pin.t14 0.41
R365 pin.n70 pin.t15 0.41
R366 pin.n70 pin.t10 0.41
R367 pin.n61 pin.t214 0.41
R368 pin.n61 pin.t216 0.41
R369 pin.n60 pin.t218 0.41
R370 pin.n60 pin.t215 0.41
R371 pin.n51 pin.t179 0.41
R372 pin.n51 pin.t175 0.41
R373 pin.n50 pin.t177 0.41
R374 pin.n50 pin.t180 0.41
R375 pin.n41 pin.t62 0.41
R376 pin.n41 pin.t58 0.41
R377 pin.n40 pin.t59 0.41
R378 pin.n40 pin.t60 0.41
R379 pin.n31 pin.t200 0.41
R380 pin.n31 pin.t203 0.41
R381 pin.n30 pin.t205 0.41
R382 pin.n30 pin.t201 0.41
R383 pin.n21 pin.t171 0.41
R384 pin.n21 pin.t172 0.41
R385 pin.n20 pin.t174 0.41
R386 pin.n20 pin.t169 0.41
R387 pin.n11 pin.t64 0.41
R388 pin.n11 pin.t66 0.41
R389 pin.n10 pin.t67 0.41
R390 pin.n10 pin.t65 0.41
R391 pin.n1 pin.t196 0.41
R392 pin.n1 pin.t199 0.41
R393 pin.n0 pin.t195 0.41
R394 pin.n0 pin.t197 0.41
R395 pin.n113 pin.n112 0.230427
R396 pin.n126 pin.n125 0.230427
R397 pin.n139 pin.n138 0.230427
R398 pin.n152 pin.n151 0.230427
R399 pin.n165 pin.n164 0.230427
R400 pin.n178 pin.n177 0.230427
R401 pin.n191 pin.n190 0.230427
R402 pin.n204 pin.n203 0.230427
R403 pin.n217 pin.n216 0.230427
R404 pin.n109 pin.n108 0.22977
R405 pin.n122 pin.n121 0.22977
R406 pin.n135 pin.n134 0.22977
R407 pin.n148 pin.n147 0.22977
R408 pin.n161 pin.n160 0.22977
R409 pin.n174 pin.n173 0.22977
R410 pin.n187 pin.n186 0.22977
R411 pin.n200 pin.n199 0.22977
R412 pin.n213 pin.n212 0.22977
R413 pin.n226 pin.n225 0.22977
R414 pin.n111 pin.n110 0.227799
R415 pin.n124 pin.n123 0.227799
R416 pin.n137 pin.n136 0.227799
R417 pin.n150 pin.n149 0.227799
R418 pin.n163 pin.n162 0.227799
R419 pin.n176 pin.n175 0.227799
R420 pin.n189 pin.n188 0.227799
R421 pin.n202 pin.n201 0.227799
R422 pin.n215 pin.n214 0.227799
R423 pin.n228 pin.n227 0.227799
R424 pin.n101 pin.n100 0.210719
R425 pin.n102 pin.n101 0.210719
R426 pin.n103 pin.n102 0.210719
R427 pin.n104 pin.n103 0.210719
R428 pin.n105 pin.n104 0.210719
R429 pin.n106 pin.n105 0.210719
R430 pin.n107 pin.n106 0.210719
R431 pin.n110 pin.n109 0.210719
R432 pin.n114 pin.n113 0.210719
R433 pin.n115 pin.n114 0.210719
R434 pin.n116 pin.n115 0.210719
R435 pin.n117 pin.n116 0.210719
R436 pin.n118 pin.n117 0.210719
R437 pin.n119 pin.n118 0.210719
R438 pin.n120 pin.n119 0.210719
R439 pin.n123 pin.n122 0.210719
R440 pin.n127 pin.n126 0.210719
R441 pin.n128 pin.n127 0.210719
R442 pin.n129 pin.n128 0.210719
R443 pin.n130 pin.n129 0.210719
R444 pin.n131 pin.n130 0.210719
R445 pin.n132 pin.n131 0.210719
R446 pin.n133 pin.n132 0.210719
R447 pin.n136 pin.n135 0.210719
R448 pin.n140 pin.n139 0.210719
R449 pin.n141 pin.n140 0.210719
R450 pin.n142 pin.n141 0.210719
R451 pin.n143 pin.n142 0.210719
R452 pin.n144 pin.n143 0.210719
R453 pin.n145 pin.n144 0.210719
R454 pin.n146 pin.n145 0.210719
R455 pin.n149 pin.n148 0.210719
R456 pin.n153 pin.n152 0.210719
R457 pin.n154 pin.n153 0.210719
R458 pin.n155 pin.n154 0.210719
R459 pin.n156 pin.n155 0.210719
R460 pin.n157 pin.n156 0.210719
R461 pin.n158 pin.n157 0.210719
R462 pin.n159 pin.n158 0.210719
R463 pin.n162 pin.n161 0.210719
R464 pin.n166 pin.n165 0.210719
R465 pin.n167 pin.n166 0.210719
R466 pin.n168 pin.n167 0.210719
R467 pin.n169 pin.n168 0.210719
R468 pin.n170 pin.n169 0.210719
R469 pin.n171 pin.n170 0.210719
R470 pin.n172 pin.n171 0.210719
R471 pin.n175 pin.n174 0.210719
R472 pin.n179 pin.n178 0.210719
R473 pin.n180 pin.n179 0.210719
R474 pin.n181 pin.n180 0.210719
R475 pin.n182 pin.n181 0.210719
R476 pin.n183 pin.n182 0.210719
R477 pin.n184 pin.n183 0.210719
R478 pin.n185 pin.n184 0.210719
R479 pin.n188 pin.n187 0.210719
R480 pin.n192 pin.n191 0.210719
R481 pin.n193 pin.n192 0.210719
R482 pin.n194 pin.n193 0.210719
R483 pin.n195 pin.n194 0.210719
R484 pin.n196 pin.n195 0.210719
R485 pin.n197 pin.n196 0.210719
R486 pin.n198 pin.n197 0.210719
R487 pin.n201 pin.n200 0.210719
R488 pin.n205 pin.n204 0.210719
R489 pin.n206 pin.n205 0.210719
R490 pin.n207 pin.n206 0.210719
R491 pin.n208 pin.n207 0.210719
R492 pin.n209 pin.n208 0.210719
R493 pin.n210 pin.n209 0.210719
R494 pin.n211 pin.n210 0.210719
R495 pin.n214 pin.n213 0.210719
R496 pin.n218 pin.n217 0.210719
R497 pin.n219 pin.n218 0.210719
R498 pin.n220 pin.n219 0.210719
R499 pin.n221 pin.n220 0.210719
R500 pin.n222 pin.n221 0.210719
R501 pin.n223 pin.n222 0.210719
R502 pin.n224 pin.n223 0.210719
R503 pin.n227 pin.n226 0.210719
R504 BUS[5].n5 BUS[5].t11 15.5918
R505 BUS[5].n2 BUS[5].n0 15.3751
R506 BUS[5].n8 BUS[5].n6 15.2168
R507 BUS[5].n2 BUS[5].n1 15.0151
R508 BUS[5].n4 BUS[5].n3 15.0151
R509 BUS[5].n20 BUS[5].n19 14.8568
R510 BUS[5].n18 BUS[5].n17 14.8568
R511 BUS[5].n16 BUS[5].n15 14.8568
R512 BUS[5].n14 BUS[5].n13 14.8568
R513 BUS[5].n12 BUS[5].n11 14.8568
R514 BUS[5].n10 BUS[5].n9 14.8568
R515 BUS[5].n8 BUS[5].n7 14.8568
R516 BUS[5].n21 BUS[5] 0.921051
R517 BUS[5].n5 BUS[5].n4 0.8465
R518 BUS[5].n19 BUS[5].t1 0.4555
R519 BUS[5].n19 BUS[5].t9 0.4555
R520 BUS[5].n17 BUS[5].t13 0.4555
R521 BUS[5].n17 BUS[5].t10 0.4555
R522 BUS[5].n15 BUS[5].t3 0.4555
R523 BUS[5].n15 BUS[5].t6 0.4555
R524 BUS[5].n13 BUS[5].t5 0.4555
R525 BUS[5].n13 BUS[5].t12 0.4555
R526 BUS[5].n11 BUS[5].t0 0.4555
R527 BUS[5].n11 BUS[5].t2 0.4555
R528 BUS[5].n9 BUS[5].t8 0.4555
R529 BUS[5].n9 BUS[5].t15 0.4555
R530 BUS[5].n7 BUS[5].t14 0.4555
R531 BUS[5].n7 BUS[5].t16 0.4555
R532 BUS[5].n6 BUS[5].t4 0.4555
R533 BUS[5].n6 BUS[5].t7 0.4555
R534 BUS[5].n0 BUS[5].t22 0.41
R535 BUS[5].n0 BUS[5].t17 0.41
R536 BUS[5].n1 BUS[5].t19 0.41
R537 BUS[5].n1 BUS[5].t21 0.41
R538 BUS[5].n3 BUS[5].t20 0.41
R539 BUS[5].n3 BUS[5].t18 0.41
R540 BUS[5].n4 BUS[5].n2 0.3605
R541 BUS[5].n10 BUS[5].n8 0.3605
R542 BUS[5].n12 BUS[5].n10 0.3605
R543 BUS[5].n14 BUS[5].n12 0.3605
R544 BUS[5].n16 BUS[5].n14 0.3605
R545 BUS[5].n18 BUS[5].n16 0.3605
R546 BUS[5].n20 BUS[5].n18 0.3605
R547 BUS[5].n21 BUS[5].n5 0.14225
R548 BUS[5].n21 BUS[5].n20 0.111875
R549 BUS[5] BUS[5].n21 0.044437
R550 vdd.t218 vdd.t216 667.707
R551 vdd.t100 vdd.t102 667.707
R552 vdd.t385 vdd.t383 667.707
R553 vdd.t198 vdd.t196 667.707
R554 vdd.t204 vdd.t206 667.707
R555 vdd.t15 vdd.t17 667.707
R556 vdd.t397 vdd.t399 667.707
R557 vdd.t163 vdd.t165 667.707
R558 vdd.t480 vdd.t478 667.707
R559 vdd.t377 vdd.t375 667.707
R560 vdd.t363 vdd.t361 667.707
R561 vdd.t425 vdd.t423 667.707
R562 vdd.t55 vdd.t53 667.707
R563 vdd.t89 vdd.t91 667.707
R564 vdd.t123 vdd.t121 667.707
R565 vdd.t30 vdd.t28 667.707
R566 vdd.t176 vdd.t174 667.707
R567 vdd.t238 vdd.t240 667.707
R568 vdd.t271 vdd.t269 667.707
R569 vdd.t127 vdd.t129 667.707
R570 vdd.t500 vdd.t433 574.104
R571 vdd.t9 vdd.t474 574.104
R572 vdd.t200 vdd.t278 574.104
R573 vdd.t440 vdd.t143 574.104
R574 vdd.t181 vdd.t435 574.104
R575 vdd.t387 vdd.t147 574.104
R576 vdd.t178 vdd.t405 574.104
R577 vdd.t293 vdd.t333 574.104
R578 vdd.t401 vdd.t189 574.104
R579 vdd.t154 vdd.t138 574.104
R580 vdd.t208 vdd.t131 574.104
R581 vdd.t265 vdd.t416 574.104
R582 vdd.t170 vdd.t259 574.104
R583 vdd.t511 vdd.t159 574.104
R584 vdd.t470 vdd.t329 574.104
R585 vdd.t38 vdd.t59 574.104
R586 vdd.t51 vdd.t420 574.104
R587 vdd.t446 vdd.t368 574.104
R588 vdd.t450 vdd.t98 574.104
R589 vdd.t516 vdd.t7 574.104
R590 vdd.n68 vdd.t410 569.532
R591 vdd.n61 vdd.t167 564.744
R592 vdd.n54 vdd.t427 564.744
R593 vdd.n47 vdd.t505 564.744
R594 vdd.n40 vdd.t381 564.744
R595 vdd.n33 vdd.t125 564.744
R596 vdd.n26 vdd.t111 564.744
R597 vdd.n19 vdd.t119 564.744
R598 vdd.n12 vdd.t64 564.744
R599 vdd.n5 vdd.t172 564.744
R600 vdd.n208 vdd.t106 530.606
R601 vdd.n211 vdd.t489 530.606
R602 vdd.n214 vdd.t26 530.606
R603 vdd.n217 vdd.t498 530.606
R604 vdd.n220 vdd.t392 530.606
R605 vdd.n223 vdd.t150 530.606
R606 vdd.n226 vdd.t484 530.606
R607 vdd.n229 vdd.t379 530.606
R608 vdd.n232 vdd.t152 530.606
R609 vdd.n235 vdd.t454 530.606
R610 vdd.n62 vdd.n61 474.26
R611 vdd.n55 vdd.n54 474.26
R612 vdd.n48 vdd.n47 474.26
R613 vdd.n41 vdd.n40 474.26
R614 vdd.n34 vdd.n33 474.26
R615 vdd.n27 vdd.n26 474.26
R616 vdd.n20 vdd.n19 474.26
R617 vdd.n13 vdd.n12 474.26
R618 vdd.n6 vdd.n5 474.26
R619 vdd.n65 vdd.t100 471.139
R620 vdd.n58 vdd.t198 471.139
R621 vdd.n51 vdd.t15 471.139
R622 vdd.n44 vdd.t163 471.139
R623 vdd.n37 vdd.t377 471.139
R624 vdd.n30 vdd.t425 471.139
R625 vdd.n23 vdd.t89 471.139
R626 vdd.n16 vdd.t30 471.139
R627 vdd.n9 vdd.t238 471.139
R628 vdd.n2 vdd.t127 471.139
R629 vdd vdd.t218 410.296
R630 vdd vdd.t385 410.296
R631 vdd vdd.t204 410.296
R632 vdd vdd.t397 410.296
R633 vdd vdd.t480 410.296
R634 vdd vdd.t363 410.296
R635 vdd vdd.t55 410.296
R636 vdd vdd.t123 410.296
R637 vdd vdd.t176 410.296
R638 vdd vdd.t271 410.296
R639 vdd.t433 vdd.t36 405.616
R640 vdd.t474 vdd.t302 405.616
R641 vdd.t278 vdd.t343 405.616
R642 vdd.t143 vdd.t444 405.616
R643 vdd.t435 vdd.t32 405.616
R644 vdd.t147 vdd.t526 405.616
R645 vdd.t405 vdd.t145 405.616
R646 vdd.t333 vdd.t300 405.616
R647 vdd.t189 vdd.t345 405.616
R648 vdd.t138 vdd.t256 405.616
R649 vdd.t131 vdd.t289 405.616
R650 vdd.t416 vdd.t66 405.616
R651 vdd.t259 vdd.t34 405.616
R652 vdd.t159 vdd.t68 405.616
R653 vdd.t329 vdd.t252 405.616
R654 vdd.t59 vdd.t494 405.616
R655 vdd.t420 vdd.t254 405.616
R656 vdd.t368 vdd.t528 405.616
R657 vdd.t98 vdd.t242 405.616
R658 vdd.t7 vdd.t496 405.616
R659 vdd vdd.t461 390.017
R660 vdd vdd.t463 390.017
R661 vdd vdd.t466 390.017
R662 vdd vdd.t482 390.017
R663 vdd vdd.t19 390.017
R664 vdd vdd.t457 390.017
R665 vdd vdd.t468 390.017
R666 vdd vdd.t476 390.017
R667 vdd vdd.t459 390.017
R668 vdd vdd.t21 390.017
R669 vdd.t523 vdd.t456 374.416
R670 vdd.t210 vdd.t472 374.416
R671 vdd.t57 vdd.t403 374.416
R672 vdd.t70 vdd.t141 374.416
R673 vdd.t306 vdd.t486 374.416
R674 vdd.t250 vdd.t63 374.416
R675 vdd.t331 vdd.t23 374.416
R676 vdd.t371 vdd.t169 374.416
R677 vdd.t93 vdd.t429 374.416
R678 vdd.t336 vdd.t338 374.416
R679 vdd.t95 vdd.t62 374.416
R680 vdd.t491 vdd.t391 374.416
R681 vdd.t161 vdd.t180 374.416
R682 vdd.t502 vdd.t110 374.416
R683 vdd.t134 vdd.t137 374.416
R684 vdd.t487 vdd.t515 374.416
R685 vdd.t191 vdd.t212 374.416
R686 vdd.t221 vdd.t136 374.416
R687 vdd.t412 vdd.t215 374.416
R688 vdd.t452 vdd.t465 374.416
R689 vdd.t461 vdd.t340 318.253
R690 vdd.t216 vdd.t523 318.253
R691 vdd.t456 vdd.t432 318.253
R692 vdd.t102 vdd.t210 318.253
R693 vdd.t472 vdd.t473 318.253
R694 vdd.t463 vdd.t11 318.253
R695 vdd.t383 vdd.t57 318.253
R696 vdd.t403 vdd.t280 318.253
R697 vdd.t196 vdd.t70 318.253
R698 vdd.t141 vdd.t142 318.253
R699 vdd.t466 vdd.t442 318.253
R700 vdd.t206 vdd.t306 318.253
R701 vdd.t486 vdd.t437 318.253
R702 vdd.t17 vdd.t250 318.253
R703 vdd.t63 vdd.t149 318.253
R704 vdd.t482 vdd.t389 318.253
R705 vdd.t399 vdd.t331 318.253
R706 vdd.t23 vdd.t404 318.253
R707 vdd.t165 vdd.t371 318.253
R708 vdd.t169 vdd.t335 318.253
R709 vdd.t19 vdd.t291 318.253
R710 vdd.t478 vdd.t93 318.253
R711 vdd.t429 vdd.t188 318.253
R712 vdd.t375 vdd.t336 318.253
R713 vdd.t338 vdd.t140 318.253
R714 vdd.t457 vdd.t156 318.253
R715 vdd.t361 vdd.t95 318.253
R716 vdd.t62 vdd.t133 318.253
R717 vdd.t423 vdd.t491 318.253
R718 vdd.t391 vdd.t418 318.253
R719 vdd.t468 vdd.t267 318.253
R720 vdd.t53 vdd.t161 318.253
R721 vdd.t180 vdd.t258 318.253
R722 vdd.t91 vdd.t502 318.253
R723 vdd.t110 vdd.t158 318.253
R724 vdd.t476 vdd.t509 318.253
R725 vdd.t121 vdd.t134 318.253
R726 vdd.t137 vdd.t328 318.253
R727 vdd.t28 vdd.t487 318.253
R728 vdd.t515 vdd.t61 318.253
R729 vdd.t459 vdd.t40 318.253
R730 vdd.t174 vdd.t191 318.253
R731 vdd.t212 vdd.t419 318.253
R732 vdd.t240 vdd.t221 318.253
R733 vdd.t136 vdd.t370 318.253
R734 vdd.t21 vdd.t448 318.253
R735 vdd.t269 vdd.t412 318.253
R736 vdd.t215 vdd.t97 318.253
R737 vdd.t129 vdd.t452 318.253
R738 vdd.t465 vdd.t6 318.253
R739 vdd.n206 vdd 293.171
R740 vdd vdd.n65 288.613
R741 vdd vdd.n62 288.613
R742 vdd vdd.n58 288.613
R743 vdd vdd.n55 288.613
R744 vdd vdd.n51 288.613
R745 vdd vdd.n48 288.613
R746 vdd vdd.n44 288.613
R747 vdd vdd.n41 288.613
R748 vdd vdd.n37 288.613
R749 vdd vdd.n34 288.613
R750 vdd vdd.n30 288.613
R751 vdd vdd.n27 288.613
R752 vdd vdd.n23 288.613
R753 vdd vdd.n20 288.613
R754 vdd vdd.n16 288.613
R755 vdd vdd.n13 288.613
R756 vdd vdd.n9 288.613
R757 vdd vdd.n6 288.613
R758 vdd vdd.n2 288.613
R759 vdd.n207 vdd.t224 243.641
R760 vdd.n209 vdd.t358 242.278
R761 vdd.n212 vdd.t115 242.278
R762 vdd.n215 vdd.t304 242.278
R763 vdd.n218 vdd.t493 242.278
R764 vdd.n221 vdd.t76 242.278
R765 vdd.n224 vdd.t373 242.278
R766 vdd.n227 vdd.t248 242.278
R767 vdd.n230 vdd.t117 242.278
R768 vdd.n233 vdd.t44 242.278
R769 vdd.t432 vdd.t500 230.889
R770 vdd.t473 vdd.t9 230.889
R771 vdd.t280 vdd.t200 230.889
R772 vdd.t142 vdd.t440 230.889
R773 vdd.t437 vdd.t181 230.889
R774 vdd.t149 vdd.t387 230.889
R775 vdd.t404 vdd.t178 230.889
R776 vdd.t335 vdd.t293 230.889
R777 vdd.t188 vdd.t401 230.889
R778 vdd.t140 vdd.t154 230.889
R779 vdd.t133 vdd.t208 230.889
R780 vdd.t418 vdd.t265 230.889
R781 vdd.t258 vdd.t170 230.889
R782 vdd.t158 vdd.t511 230.889
R783 vdd.t328 vdd.t470 230.889
R784 vdd.t61 vdd.t38 230.889
R785 vdd.t419 vdd.t51 230.889
R786 vdd.t370 vdd.t446 230.889
R787 vdd.t97 vdd.t450 230.889
R788 vdd.t6 vdd.t516 230.889
R789 vdd.t410 vdd 195.008
R790 vdd.t36 vdd 195.008
R791 vdd.t302 vdd 195.008
R792 vdd.t167 vdd 195.008
R793 vdd.t343 vdd 195.008
R794 vdd.t444 vdd 195.008
R795 vdd.t427 vdd 195.008
R796 vdd.t32 vdd 195.008
R797 vdd.t526 vdd 195.008
R798 vdd.t505 vdd 195.008
R799 vdd.t145 vdd 195.008
R800 vdd.t300 vdd 195.008
R801 vdd.t381 vdd 195.008
R802 vdd.t345 vdd 195.008
R803 vdd.t256 vdd 195.008
R804 vdd.t125 vdd 195.008
R805 vdd.t289 vdd 195.008
R806 vdd.t66 vdd 195.008
R807 vdd.t111 vdd 195.008
R808 vdd.t34 vdd 195.008
R809 vdd.t68 vdd 195.008
R810 vdd.t119 vdd 195.008
R811 vdd.t252 vdd 195.008
R812 vdd.t494 vdd 195.008
R813 vdd.t64 vdd 195.008
R814 vdd.t254 vdd 195.008
R815 vdd.t528 vdd 195.008
R816 vdd.t172 vdd 195.008
R817 vdd.t242 vdd 195.008
R818 vdd.t496 vdd 195.008
R819 vdd.t340 vdd 165.368
R820 vdd.t11 vdd 165.368
R821 vdd.t442 vdd 165.368
R822 vdd.t389 vdd 165.368
R823 vdd.t291 vdd 165.368
R824 vdd.t156 vdd 165.368
R825 vdd.t267 vdd 165.368
R826 vdd.t509 vdd 165.368
R827 vdd.t40 vdd 165.368
R828 vdd.t448 vdd 165.368
R829 vdd.t106 vdd 158.228
R830 vdd.t489 vdd 158.228
R831 vdd.t26 vdd 158.228
R832 vdd.t498 vdd 158.228
R833 vdd.t392 vdd 158.228
R834 vdd.t150 vdd 158.228
R835 vdd.t484 vdd 158.228
R836 vdd.t379 vdd 158.228
R837 vdd.t152 vdd 158.228
R838 vdd.t454 vdd 158.228
R839 vdd.t224 vdd.t277 148.7
R840 vdd.t277 vdd.t355 148.7
R841 vdd.t355 vdd.t359 148.7
R842 vdd.t359 vdd.t319 148.7
R843 vdd.t319 vdd.t354 148.7
R844 vdd.t354 vdd.t422 148.7
R845 vdd.t422 vdd.t318 148.7
R846 vdd.t318 vdd.t276 148.7
R847 vdd.t276 vdd.t213 148.7
R848 vdd.t213 vdd.t223 148.7
R849 vdd.t223 vdd.t367 148.7
R850 vdd.t367 vdd.t327 148.7
R851 vdd.t327 vdd.t326 148.7
R852 vdd.t326 vdd.t305 148.7
R853 vdd.t305 vdd.t360 148.7
R854 vdd.t360 vdd.t214 148.7
R855 vdd.t358 vdd.t202 148.7
R856 vdd.t202 vdd.t298 148.7
R857 vdd.t298 vdd.t357 148.7
R858 vdd.t357 vdd.t295 148.7
R859 vdd.t295 vdd.t339 148.7
R860 vdd.t339 vdd.t314 148.7
R861 vdd.t314 vdd.t353 148.7
R862 vdd.t353 vdd.t414 148.7
R863 vdd.t414 vdd.t508 148.7
R864 vdd.t508 vdd.t352 148.7
R865 vdd.t352 vdd.t203 148.7
R866 vdd.t203 vdd.t299 148.7
R867 vdd.t299 vdd.t273 148.7
R868 vdd.t273 vdd.t365 148.7
R869 vdd.t365 vdd.t415 148.7
R870 vdd.t415 vdd.t315 148.7
R871 vdd.t115 vdd.t13 148.7
R872 vdd.t13 vdd.t407 148.7
R873 vdd.t407 vdd.t263 148.7
R874 vdd.t263 vdd.t525 148.7
R875 vdd.t525 vdd.t281 148.7
R876 vdd.t281 vdd.t409 148.7
R877 vdd.t409 vdd.t283 148.7
R878 vdd.t283 vdd.t14 148.7
R879 vdd.t14 vdd.t408 148.7
R880 vdd.t408 vdd.t116 148.7
R881 vdd.t116 vdd.t262 148.7
R882 vdd.t262 vdd.t187 148.7
R883 vdd.t187 vdd.t186 148.7
R884 vdd.t186 vdd.t261 148.7
R885 vdd.t261 vdd.t282 148.7
R886 vdd.t282 vdd.t185 148.7
R887 vdd.t304 vdd.t366 148.7
R888 vdd.t366 vdd.t324 148.7
R889 vdd.t324 vdd.t232 148.7
R890 vdd.t232 vdd.t317 148.7
R891 vdd.t317 vdd.t296 148.7
R892 vdd.t296 vdd.t347 148.7
R893 vdd.t347 vdd.t316 148.7
R894 vdd.t316 vdd.t348 148.7
R895 vdd.t348 vdd.t342 148.7
R896 vdd.t342 vdd.t514 148.7
R897 vdd.t514 vdd.t275 148.7
R898 vdd.t275 vdd.t504 148.7
R899 vdd.t504 vdd.t513 148.7
R900 vdd.t513 vdd.t274 148.7
R901 vdd.t274 vdd.t297 148.7
R902 vdd.t297 vdd.t325 148.7
R903 vdd.t493 vdd.t244 148.7
R904 vdd.t244 vdd.t246 148.7
R905 vdd.t246 vdd.t48 148.7
R906 vdd.t48 vdd.t395 148.7
R907 vdd.t395 vdd.t245 148.7
R908 vdd.t245 vdd.t351 148.7
R909 vdd.t351 vdd.t349 148.7
R910 vdd.t349 vdd.t284 148.7
R911 vdd.t284 vdd.t236 148.7
R912 vdd.t236 vdd.t50 148.7
R913 vdd.t50 vdd.t396 148.7
R914 vdd.t396 vdd.t394 148.7
R915 vdd.t394 vdd.t49 148.7
R916 vdd.t49 vdd.t350 148.7
R917 vdd.t350 vdd.t285 148.7
R918 vdd.t285 vdd.t237 148.7
R919 vdd.t76 vdd.t79 148.7
R920 vdd.t79 vdd.t86 148.7
R921 vdd.t86 vdd.t88 148.7
R922 vdd.t88 vdd.t80 148.7
R923 vdd.t80 vdd.t87 148.7
R924 vdd.t87 vdd.t72 148.7
R925 vdd.t72 vdd.t74 148.7
R926 vdd.t74 vdd.t77 148.7
R927 vdd.t77 vdd.t84 148.7
R928 vdd.t84 vdd.t75 148.7
R929 vdd.t75 vdd.t78 148.7
R930 vdd.t78 vdd.t85 148.7
R931 vdd.t85 vdd.t82 148.7
R932 vdd.t82 vdd.t73 148.7
R933 vdd.t73 vdd.t81 148.7
R934 vdd.t81 vdd.t83 148.7
R935 vdd.t373 vdd.t320 148.7
R936 vdd.t320 vdd.t310 148.7
R937 vdd.t310 vdd.t313 148.7
R938 vdd.t313 vdd.t183 148.7
R939 vdd.t183 vdd.t439 148.7
R940 vdd.t439 vdd.t356 148.7
R941 vdd.t356 vdd.t321 148.7
R942 vdd.t321 vdd.t438 148.7
R943 vdd.t438 vdd.t311 148.7
R944 vdd.t311 vdd.t374 148.7
R945 vdd.t374 vdd.t312 148.7
R946 vdd.t312 vdd.t309 148.7
R947 vdd.t309 vdd.t323 148.7
R948 vdd.t323 vdd.t264 148.7
R949 vdd.t264 vdd.t308 148.7
R950 vdd.t308 vdd.t322 148.7
R951 vdd.t248 vdd.t45 148.7
R952 vdd.t45 vdd.t249 148.7
R953 vdd.t249 vdd.t247 148.7
R954 vdd.t247 vdd.t231 148.7
R955 vdd.t231 vdd.t47 148.7
R956 vdd.t47 vdd.t234 148.7
R957 vdd.t234 vdd.t230 148.7
R958 vdd.t230 vdd.t46 148.7
R959 vdd.t46 vdd.t233 148.7
R960 vdd.t233 vdd.t184 148.7
R961 vdd.t184 vdd.t431 148.7
R962 vdd.t431 vdd.t113 148.7
R963 vdd.t113 vdd.t235 148.7
R964 vdd.t235 vdd.t430 148.7
R965 vdd.t430 vdd.t229 148.7
R966 vdd.t229 vdd.t114 148.7
R967 vdd.t117 vdd.t3 148.7
R968 vdd.t3 vdd.t195 148.7
R969 vdd.t195 vdd.t25 148.7
R970 vdd.t25 vdd.t104 148.7
R971 vdd.t104 vdd.t507 148.7
R972 vdd.t507 vdd.t220 148.7
R973 vdd.t220 vdd.t118 148.7
R974 vdd.t118 vdd.t4 148.7
R975 vdd.t4 vdd.t1 148.7
R976 vdd.t1 vdd.t194 148.7
R977 vdd.t194 vdd.t24 148.7
R978 vdd.t24 vdd.t0 148.7
R979 vdd.t0 vdd.t193 148.7
R980 vdd.t193 vdd.t105 148.7
R981 vdd.t105 vdd.t5 148.7
R982 vdd.t5 vdd.t2 148.7
R983 vdd.t44 vdd.t228 148.7
R984 vdd.t228 vdd.t288 148.7
R985 vdd.t288 vdd.t43 148.7
R986 vdd.t43 vdd.t42 148.7
R987 vdd.t42 vdd.t287 148.7
R988 vdd.t287 vdd.t521 148.7
R989 vdd.t521 vdd.t519 148.7
R990 vdd.t519 vdd.t226 148.7
R991 vdd.t226 vdd.t109 148.7
R992 vdd.t109 vdd.t518 148.7
R993 vdd.t518 vdd.t225 148.7
R994 vdd.t225 vdd.t108 148.7
R995 vdd.t108 vdd.t286 148.7
R996 vdd.t286 vdd.t520 148.7
R997 vdd.t520 vdd.t227 148.7
R998 vdd.t227 vdd.t522 148.7
R999 vdd.n195 vdd.t22 15.5636
R1000 vdd.n181 vdd.t460 15.5636
R1001 vdd.n167 vdd.t477 15.5636
R1002 vdd.n153 vdd.t469 15.5636
R1003 vdd.n139 vdd.t458 15.5636
R1004 vdd.n125 vdd.t20 15.5636
R1005 vdd.n111 vdd.t483 15.5636
R1006 vdd.n97 vdd.t467 15.5636
R1007 vdd.n83 vdd.t464 15.5636
R1008 vdd.n69 vdd.t462 15.5636
R1009 vdd.n204 vdd.t517 4.77854
R1010 vdd.n199 vdd.t451 4.77854
R1011 vdd.n190 vdd.t447 4.77854
R1012 vdd.n185 vdd.t52 4.77854
R1013 vdd.n176 vdd.t39 4.77854
R1014 vdd.n171 vdd.t471 4.77854
R1015 vdd.n162 vdd.t512 4.77854
R1016 vdd.n157 vdd.t171 4.77854
R1017 vdd.n148 vdd.t266 4.77854
R1018 vdd.n143 vdd.t209 4.77854
R1019 vdd.n134 vdd.t155 4.77854
R1020 vdd.n129 vdd.t402 4.77854
R1021 vdd.n120 vdd.t294 4.77854
R1022 vdd.n115 vdd.t179 4.77854
R1023 vdd.n106 vdd.t388 4.77854
R1024 vdd.n101 vdd.t182 4.77854
R1025 vdd.n92 vdd.t441 4.77854
R1026 vdd.n87 vdd.t201 4.77854
R1027 vdd.n78 vdd.t10 4.77854
R1028 vdd.n73 vdd.t501 4.77854
R1029 vdd.n201 vdd.n2 4.55932
R1030 vdd.n193 vdd.n5 4.55932
R1031 vdd.n192 vdd.n6 4.55932
R1032 vdd.n187 vdd.n9 4.55932
R1033 vdd.n179 vdd.n12 4.55932
R1034 vdd.n178 vdd.n13 4.55932
R1035 vdd.n173 vdd.n16 4.55932
R1036 vdd.n165 vdd.n19 4.55932
R1037 vdd.n164 vdd.n20 4.55932
R1038 vdd.n159 vdd.n23 4.55932
R1039 vdd.n151 vdd.n26 4.55932
R1040 vdd.n150 vdd.n27 4.55932
R1041 vdd.n145 vdd.n30 4.55932
R1042 vdd.n137 vdd.n33 4.55932
R1043 vdd.n136 vdd.n34 4.55932
R1044 vdd.n131 vdd.n37 4.55932
R1045 vdd.n123 vdd.n40 4.55932
R1046 vdd.n122 vdd.n41 4.55932
R1047 vdd.n117 vdd.n44 4.55932
R1048 vdd.n109 vdd.n47 4.55932
R1049 vdd.n108 vdd.n48 4.55932
R1050 vdd.n103 vdd.n51 4.55932
R1051 vdd.n95 vdd.n54 4.55932
R1052 vdd.n94 vdd.n55 4.55932
R1053 vdd.n89 vdd.n58 4.55932
R1054 vdd.n81 vdd.n61 4.55932
R1055 vdd.n80 vdd.n62 4.55932
R1056 vdd.n75 vdd.n65 4.55932
R1057 vdd.n202 vdd.t128 3.95308
R1058 vdd.n197 vdd.t272 3.95308
R1059 vdd.n188 vdd.t239 3.95308
R1060 vdd.n183 vdd.t177 3.95308
R1061 vdd.n174 vdd.t31 3.95308
R1062 vdd.n169 vdd.t124 3.95308
R1063 vdd.n160 vdd.t90 3.95308
R1064 vdd.n155 vdd.t56 3.95308
R1065 vdd.n146 vdd.t426 3.95308
R1066 vdd.n141 vdd.t364 3.95308
R1067 vdd.n132 vdd.t378 3.95308
R1068 vdd.n127 vdd.t481 3.95308
R1069 vdd.n118 vdd.t164 3.95308
R1070 vdd.n113 vdd.t398 3.95308
R1071 vdd.n104 vdd.t16 3.95308
R1072 vdd.n99 vdd.t205 3.95308
R1073 vdd.n90 vdd.t199 3.95308
R1074 vdd.n85 vdd.t386 3.95308
R1075 vdd.n76 vdd.t101 3.95308
R1076 vdd.n71 vdd.t219 3.95308
R1077 vdd.n196 vdd.t449 3.90058
R1078 vdd.n182 vdd.t41 3.90058
R1079 vdd.n168 vdd.t510 3.90058
R1080 vdd.n154 vdd.t268 3.90058
R1081 vdd.n140 vdd.t157 3.90058
R1082 vdd.n126 vdd.t292 3.90058
R1083 vdd.n112 vdd.t390 3.90058
R1084 vdd.n98 vdd.t443 3.90058
R1085 vdd.n84 vdd.t12 3.90058
R1086 vdd.n70 vdd.t341 3.90058
R1087 vdd.n207 vdd.t107 3.84351
R1088 vdd.n210 vdd.t490 3.84351
R1089 vdd.n213 vdd.t27 3.84351
R1090 vdd.n216 vdd.t499 3.84351
R1091 vdd.n219 vdd.t393 3.84351
R1092 vdd.n222 vdd.t151 3.84351
R1093 vdd.n225 vdd.t485 3.84351
R1094 vdd.n228 vdd.t380 3.84351
R1095 vdd.n231 vdd.t153 3.84351
R1096 vdd.n234 vdd.t455 3.84351
R1097 vdd.n194 vdd.t173 3.84351
R1098 vdd.n180 vdd.t65 3.84351
R1099 vdd.n166 vdd.t120 3.84351
R1100 vdd.n152 vdd.t112 3.84351
R1101 vdd.n138 vdd.t126 3.84351
R1102 vdd.n124 vdd.t382 3.84351
R1103 vdd.n110 vdd.t506 3.84351
R1104 vdd.n96 vdd.t428 3.84351
R1105 vdd.n82 vdd.t168 3.84351
R1106 vdd.n68 vdd.t411 3.84351
R1107 vdd.n0 vdd.t8 3.7805
R1108 vdd.n3 vdd.t99 3.7805
R1109 vdd.n7 vdd.t369 3.7805
R1110 vdd.n10 vdd.t421 3.7805
R1111 vdd.n14 vdd.t60 3.7805
R1112 vdd.n17 vdd.t330 3.7805
R1113 vdd.n21 vdd.t160 3.7805
R1114 vdd.n24 vdd.t260 3.7805
R1115 vdd.n28 vdd.t417 3.7805
R1116 vdd.n31 vdd.t132 3.7805
R1117 vdd.n35 vdd.t139 3.7805
R1118 vdd.n38 vdd.t190 3.7805
R1119 vdd.n42 vdd.t334 3.7805
R1120 vdd.n45 vdd.t406 3.7805
R1121 vdd.n49 vdd.t148 3.7805
R1122 vdd.n52 vdd.t436 3.7805
R1123 vdd.n56 vdd.t144 3.7805
R1124 vdd.n59 vdd.t279 3.7805
R1125 vdd.n63 vdd.t475 3.7805
R1126 vdd.n66 vdd.t434 3.7805
R1127 vdd.n205 vdd.n0 2.95854
R1128 vdd.n203 vdd.n1 2.95854
R1129 vdd.n200 vdd.n3 2.95854
R1130 vdd.n198 vdd.n4 2.95854
R1131 vdd.n191 vdd.n7 2.95854
R1132 vdd.n189 vdd.n8 2.95854
R1133 vdd.n186 vdd.n10 2.95854
R1134 vdd.n184 vdd.n11 2.95854
R1135 vdd.n177 vdd.n14 2.95854
R1136 vdd.n175 vdd.n15 2.95854
R1137 vdd.n172 vdd.n17 2.95854
R1138 vdd.n170 vdd.n18 2.95854
R1139 vdd.n163 vdd.n21 2.95854
R1140 vdd.n161 vdd.n22 2.95854
R1141 vdd.n158 vdd.n24 2.95854
R1142 vdd.n156 vdd.n25 2.95854
R1143 vdd.n149 vdd.n28 2.95854
R1144 vdd.n147 vdd.n29 2.95854
R1145 vdd.n144 vdd.n31 2.95854
R1146 vdd.n142 vdd.n32 2.95854
R1147 vdd.n135 vdd.n35 2.95854
R1148 vdd.n133 vdd.n36 2.95854
R1149 vdd.n130 vdd.n38 2.95854
R1150 vdd.n128 vdd.n39 2.95854
R1151 vdd.n121 vdd.n42 2.95854
R1152 vdd.n119 vdd.n43 2.95854
R1153 vdd.n116 vdd.n45 2.95854
R1154 vdd.n114 vdd.n46 2.95854
R1155 vdd.n107 vdd.n49 2.95854
R1156 vdd.n105 vdd.n50 2.95854
R1157 vdd.n102 vdd.n52 2.95854
R1158 vdd.n100 vdd.n53 2.95854
R1159 vdd.n93 vdd.n56 2.95854
R1160 vdd.n91 vdd.n57 2.95854
R1161 vdd.n88 vdd.n59 2.95854
R1162 vdd.n86 vdd.n60 2.95854
R1163 vdd.n79 vdd.n63 2.95854
R1164 vdd.n77 vdd.n64 2.95854
R1165 vdd.n74 vdd.n66 2.95854
R1166 vdd.n72 vdd.n67 2.95854
R1167 vdd.n0 vdd.t497 1.53332
R1168 vdd.n3 vdd.t243 1.53332
R1169 vdd.n7 vdd.t529 1.53332
R1170 vdd.n10 vdd.t255 1.53332
R1171 vdd.n14 vdd.t495 1.53332
R1172 vdd.n17 vdd.t253 1.53332
R1173 vdd.n21 vdd.t69 1.53332
R1174 vdd.n24 vdd.t35 1.53332
R1175 vdd.n28 vdd.t67 1.53332
R1176 vdd.n31 vdd.t290 1.53332
R1177 vdd.n35 vdd.t257 1.53332
R1178 vdd.n38 vdd.t346 1.53332
R1179 vdd.n42 vdd.t301 1.53332
R1180 vdd.n45 vdd.t146 1.53332
R1181 vdd.n49 vdd.t527 1.53332
R1182 vdd.n52 vdd.t33 1.53332
R1183 vdd.n56 vdd.t445 1.53332
R1184 vdd.n59 vdd.t344 1.53332
R1185 vdd.n63 vdd.t303 1.53332
R1186 vdd.n66 vdd.t37 1.53332
R1187 vdd.n210 vdd.n209 1.36373
R1188 vdd.n213 vdd.n212 1.36373
R1189 vdd.n216 vdd.n215 1.36373
R1190 vdd.n219 vdd.n218 1.36373
R1191 vdd.n222 vdd.n221 1.36373
R1192 vdd.n225 vdd.n224 1.36373
R1193 vdd.n228 vdd.n227 1.36373
R1194 vdd.n231 vdd.n230 1.36373
R1195 vdd.n234 vdd.n233 1.36373
R1196 vdd.n1 vdd.t130 1.31934
R1197 vdd.n1 vdd.t453 1.31934
R1198 vdd.n4 vdd.t270 1.31934
R1199 vdd.n4 vdd.t413 1.31934
R1200 vdd.n8 vdd.t241 1.31934
R1201 vdd.n8 vdd.t222 1.31934
R1202 vdd.n11 vdd.t175 1.31934
R1203 vdd.n11 vdd.t192 1.31934
R1204 vdd.n15 vdd.t29 1.31934
R1205 vdd.n15 vdd.t488 1.31934
R1206 vdd.n18 vdd.t122 1.31934
R1207 vdd.n18 vdd.t135 1.31934
R1208 vdd.n22 vdd.t92 1.31934
R1209 vdd.n22 vdd.t503 1.31934
R1210 vdd.n25 vdd.t54 1.31934
R1211 vdd.n25 vdd.t162 1.31934
R1212 vdd.n29 vdd.t424 1.31934
R1213 vdd.n29 vdd.t492 1.31934
R1214 vdd.n32 vdd.t362 1.31934
R1215 vdd.n32 vdd.t96 1.31934
R1216 vdd.n36 vdd.t376 1.31934
R1217 vdd.n36 vdd.t337 1.31934
R1218 vdd.n39 vdd.t479 1.31934
R1219 vdd.n39 vdd.t94 1.31934
R1220 vdd.n43 vdd.t166 1.31934
R1221 vdd.n43 vdd.t372 1.31934
R1222 vdd.n46 vdd.t400 1.31934
R1223 vdd.n46 vdd.t332 1.31934
R1224 vdd.n50 vdd.t18 1.31934
R1225 vdd.n50 vdd.t251 1.31934
R1226 vdd.n53 vdd.t207 1.31934
R1227 vdd.n53 vdd.t307 1.31934
R1228 vdd.n57 vdd.t197 1.31934
R1229 vdd.n57 vdd.t71 1.31934
R1230 vdd.n60 vdd.t384 1.31934
R1231 vdd.n60 vdd.t58 1.31934
R1232 vdd.n64 vdd.t103 1.31934
R1233 vdd.n64 vdd.t211 1.31934
R1234 vdd.n67 vdd.t217 1.31934
R1235 vdd.n67 vdd.t524 1.31934
R1236 vdd.n236 vdd 1.21837
R1237 vdd.n73 vdd.n72 0.3985
R1238 vdd.n78 vdd.n77 0.3985
R1239 vdd.n87 vdd.n86 0.3985
R1240 vdd.n92 vdd.n91 0.3985
R1241 vdd.n101 vdd.n100 0.3985
R1242 vdd.n106 vdd.n105 0.3985
R1243 vdd.n115 vdd.n114 0.3985
R1244 vdd.n120 vdd.n119 0.3985
R1245 vdd.n129 vdd.n128 0.3985
R1246 vdd.n134 vdd.n133 0.3985
R1247 vdd.n143 vdd.n142 0.3985
R1248 vdd.n148 vdd.n147 0.3985
R1249 vdd.n157 vdd.n156 0.3985
R1250 vdd.n162 vdd.n161 0.3985
R1251 vdd.n171 vdd.n170 0.3985
R1252 vdd.n176 vdd.n175 0.3985
R1253 vdd.n185 vdd.n184 0.3985
R1254 vdd.n190 vdd.n189 0.3985
R1255 vdd.n199 vdd.n198 0.3985
R1256 vdd.n204 vdd.n203 0.3985
R1257 vdd.n72 vdd.n71 0.3165
R1258 vdd.n77 vdd.n76 0.3165
R1259 vdd.n86 vdd.n85 0.3165
R1260 vdd.n91 vdd.n90 0.3165
R1261 vdd.n100 vdd.n99 0.3165
R1262 vdd.n105 vdd.n104 0.3165
R1263 vdd.n114 vdd.n113 0.3165
R1264 vdd.n119 vdd.n118 0.3165
R1265 vdd.n128 vdd.n127 0.3165
R1266 vdd.n133 vdd.n132 0.3165
R1267 vdd.n142 vdd.n141 0.3165
R1268 vdd.n147 vdd.n146 0.3165
R1269 vdd.n156 vdd.n155 0.3165
R1270 vdd.n161 vdd.n160 0.3165
R1271 vdd.n170 vdd.n169 0.3165
R1272 vdd.n175 vdd.n174 0.3165
R1273 vdd.n184 vdd.n183 0.3165
R1274 vdd.n189 vdd.n188 0.3165
R1275 vdd.n198 vdd.n197 0.3165
R1276 vdd.n203 vdd.n202 0.3165
R1277 vdd.n233 vdd 0.261307
R1278 vdd.n209 vdd 0.235269
R1279 vdd.n212 vdd 0.235269
R1280 vdd.n215 vdd 0.235269
R1281 vdd.n218 vdd 0.235269
R1282 vdd.n221 vdd 0.235269
R1283 vdd.n224 vdd 0.235269
R1284 vdd.n227 vdd 0.235269
R1285 vdd.n230 vdd 0.235269
R1286 vdd.n82 vdd.n81 0.2305
R1287 vdd.n96 vdd.n95 0.2305
R1288 vdd.n110 vdd.n109 0.2305
R1289 vdd.n124 vdd.n123 0.2305
R1290 vdd.n138 vdd.n137 0.2305
R1291 vdd.n152 vdd.n151 0.2305
R1292 vdd.n166 vdd.n165 0.2305
R1293 vdd.n180 vdd.n179 0.2305
R1294 vdd.n194 vdd.n193 0.2305
R1295 vdd.n74 vdd.n73 0.2125
R1296 vdd.n79 vdd.n78 0.2125
R1297 vdd.n88 vdd.n87 0.2125
R1298 vdd.n93 vdd.n92 0.2125
R1299 vdd.n102 vdd.n101 0.2125
R1300 vdd.n107 vdd.n106 0.2125
R1301 vdd.n116 vdd.n115 0.2125
R1302 vdd.n121 vdd.n120 0.2125
R1303 vdd.n130 vdd.n129 0.2125
R1304 vdd.n135 vdd.n134 0.2125
R1305 vdd.n144 vdd.n143 0.2125
R1306 vdd.n149 vdd.n148 0.2125
R1307 vdd.n158 vdd.n157 0.2125
R1308 vdd.n163 vdd.n162 0.2125
R1309 vdd.n172 vdd.n171 0.2125
R1310 vdd.n177 vdd.n176 0.2125
R1311 vdd.n186 vdd.n185 0.2125
R1312 vdd.n191 vdd.n190 0.2125
R1313 vdd.n200 vdd.n199 0.2125
R1314 vdd.n205 vdd.n204 0.2125
R1315 vdd.n75 vdd.n74 0.2085
R1316 vdd.n89 vdd.n88 0.2085
R1317 vdd.n103 vdd.n102 0.2085
R1318 vdd.n117 vdd.n116 0.2085
R1319 vdd.n131 vdd.n130 0.2085
R1320 vdd.n145 vdd.n144 0.2085
R1321 vdd.n159 vdd.n158 0.2085
R1322 vdd.n173 vdd.n172 0.2085
R1323 vdd.n187 vdd.n186 0.2085
R1324 vdd.n201 vdd.n200 0.2085
R1325 vdd.n70 vdd.n69 0.2045
R1326 vdd.n84 vdd.n83 0.2045
R1327 vdd.n98 vdd.n97 0.2045
R1328 vdd.n112 vdd.n111 0.2045
R1329 vdd.n126 vdd.n125 0.2045
R1330 vdd.n140 vdd.n139 0.2045
R1331 vdd.n154 vdd.n153 0.2045
R1332 vdd.n168 vdd.n167 0.2045
R1333 vdd.n182 vdd.n181 0.2045
R1334 vdd.n196 vdd.n195 0.2045
R1335 vdd.n80 vdd 0.1415
R1336 vdd.n94 vdd 0.1415
R1337 vdd.n108 vdd 0.1415
R1338 vdd.n122 vdd 0.1415
R1339 vdd.n136 vdd 0.1415
R1340 vdd.n150 vdd 0.1415
R1341 vdd.n164 vdd 0.1415
R1342 vdd.n178 vdd 0.1415
R1343 vdd.n192 vdd 0.1415
R1344 vdd.n206 vdd 0.1415
R1345 vdd.n76 vdd.n75 0.0985
R1346 vdd.n90 vdd.n89 0.0985
R1347 vdd.n104 vdd.n103 0.0985
R1348 vdd.n118 vdd.n117 0.0985
R1349 vdd.n132 vdd.n131 0.0985
R1350 vdd.n146 vdd.n145 0.0985
R1351 vdd.n160 vdd.n159 0.0985
R1352 vdd.n174 vdd.n173 0.0985
R1353 vdd.n188 vdd.n187 0.0985
R1354 vdd.n202 vdd.n201 0.0985
R1355 vdd vdd.n236 0.09
R1356 vdd.n69 vdd.n68 0.086
R1357 vdd.n83 vdd.n82 0.086
R1358 vdd.n97 vdd.n96 0.086
R1359 vdd.n111 vdd.n110 0.086
R1360 vdd.n125 vdd.n124 0.086
R1361 vdd.n139 vdd.n138 0.086
R1362 vdd.n153 vdd.n152 0.086
R1363 vdd.n167 vdd.n166 0.086
R1364 vdd.n181 vdd.n180 0.086
R1365 vdd.n195 vdd.n194 0.086
R1366 vdd.n71 vdd.n70 0.083
R1367 vdd.n85 vdd.n84 0.083
R1368 vdd.n99 vdd.n98 0.083
R1369 vdd.n113 vdd.n112 0.083
R1370 vdd.n127 vdd.n126 0.083
R1371 vdd.n141 vdd.n140 0.083
R1372 vdd.n155 vdd.n154 0.083
R1373 vdd.n169 vdd.n168 0.083
R1374 vdd.n183 vdd.n182 0.083
R1375 vdd.n197 vdd.n196 0.083
R1376 vdd vdd.n80 0.0775
R1377 vdd vdd.n94 0.0775
R1378 vdd vdd.n108 0.0775
R1379 vdd vdd.n122 0.0775
R1380 vdd vdd.n136 0.0775
R1381 vdd vdd.n150 0.0775
R1382 vdd vdd.n164 0.0775
R1383 vdd vdd.n178 0.0775
R1384 vdd vdd.n192 0.0775
R1385 vdd vdd.n206 0.0775
R1386 vdd.n81 vdd 0.0755
R1387 vdd.n95 vdd 0.0755
R1388 vdd.n109 vdd 0.0755
R1389 vdd.n123 vdd 0.0755
R1390 vdd.n137 vdd 0.0755
R1391 vdd.n151 vdd 0.0755
R1392 vdd.n165 vdd 0.0755
R1393 vdd.n179 vdd 0.0755
R1394 vdd.n193 vdd 0.0755
R1395 vdd.n208 vdd 0.0698976
R1396 vdd.n211 vdd 0.0698976
R1397 vdd.n214 vdd 0.0698976
R1398 vdd.n217 vdd 0.0698976
R1399 vdd.n220 vdd 0.0698976
R1400 vdd.n223 vdd 0.0698976
R1401 vdd.n226 vdd 0.0698976
R1402 vdd.n229 vdd 0.0698976
R1403 vdd.n232 vdd 0.0698976
R1404 vdd.n235 vdd 0.0698976
R1405 vdd vdd.n79 0.0675
R1406 vdd vdd.n93 0.0675
R1407 vdd vdd.n107 0.0675
R1408 vdd vdd.n121 0.0675
R1409 vdd vdd.n135 0.0675
R1410 vdd vdd.n149 0.0675
R1411 vdd vdd.n163 0.0675
R1412 vdd vdd.n177 0.0675
R1413 vdd vdd.n191 0.0675
R1414 vdd vdd.n205 0.0675
R1415 vdd vdd.n207 0.0194759
R1416 vdd vdd.n210 0.0194759
R1417 vdd vdd.n213 0.0194759
R1418 vdd vdd.n216 0.0194759
R1419 vdd vdd.n219 0.0194759
R1420 vdd vdd.n222 0.0194759
R1421 vdd vdd.n225 0.0194759
R1422 vdd vdd.n228 0.0194759
R1423 vdd vdd.n231 0.0194759
R1424 vdd vdd.n234 0.0194759
R1425 vdd.n236 vdd 0.0155
R1426 vdd vdd.n208 0.00122289
R1427 vdd vdd.n211 0.00122289
R1428 vdd vdd.n214 0.00122289
R1429 vdd vdd.n217 0.00122289
R1430 vdd vdd.n220 0.00122289
R1431 vdd vdd.n223 0.00122289
R1432 vdd vdd.n226 0.00122289
R1433 vdd vdd.n229 0.00122289
R1434 vdd vdd.n232 0.00122289
R1435 vdd vdd.n235 0.00122289
R1436 vss.n304 vss.n1 1.06994e+07
R1437 vss.n129 vss.n128 13492.4
R1438 vss.n85 vss.n83 7836.69
R1439 vss.n90 vss.n88 7736.22
R1440 vss.n95 vss.n93 7736.22
R1441 vss.n100 vss.n98 7736.22
R1442 vss.n105 vss.n103 7736.22
R1443 vss.n110 vss.n108 7736.22
R1444 vss.n115 vss.n113 7736.22
R1445 vss.n120 vss.n118 7736.22
R1446 vss.n125 vss.n123 7736.22
R1447 vss.n304 vss.n303 7598.09
R1448 vss.n90 vss.n89 3942.62
R1449 vss.n95 vss.n94 3942.62
R1450 vss.n100 vss.n99 3942.62
R1451 vss.n105 vss.n104 3942.62
R1452 vss.n110 vss.n109 3942.62
R1453 vss.n115 vss.n114 3942.62
R1454 vss.n120 vss.n119 3942.62
R1455 vss.n125 vss.n124 3942.62
R1456 vss.n85 vss.n84 3317.24
R1457 vss.n86 vss.n85 2890.76
R1458 vss.n91 vss.n90 2790.29
R1459 vss.n96 vss.n95 2790.29
R1460 vss.n101 vss.n100 2790.29
R1461 vss.n106 vss.n105 2790.29
R1462 vss.n111 vss.n110 2790.29
R1463 vss.n116 vss.n115 2790.29
R1464 vss.n121 vss.n120 2790.29
R1465 vss.n126 vss.n125 2790.29
R1466 vss.t177 vss.t179 1611.86
R1467 vss.t393 vss.t312 1611.86
R1468 vss.t269 vss.t267 1611.86
R1469 vss.t165 vss.t204 1611.86
R1470 vss.t169 vss.t167 1611.86
R1471 vss.t154 vss.t317 1611.86
R1472 vss.t284 vss.t286 1611.86
R1473 vss.t151 vss.t292 1611.86
R1474 vss.t358 vss.t356 1611.86
R1475 vss.t288 vss.t156 1611.86
R1476 vss.t244 vss.t246 1611.86
R1477 vss.t171 vss.t91 1611.86
R1478 vss.t35 vss.t37 1611.86
R1479 vss.t143 vss.t194 1611.86
R1480 vss.t80 vss.t82 1611.86
R1481 vss.t348 vss.t221 1611.86
R1482 vss.t149 vss.t147 1611.86
R1483 vss.t33 vss.t301 1611.86
R1484 vss.t200 vss.t202 1611.86
R1485 vss.t331 vss.t61 1611.86
R1486 vss.n305 vss.n304 1248.57
R1487 vss.t406 vss.t311 1138.81
R1488 vss.t312 vss.t104 1138.81
R1489 vss.t39 vss.t206 1138.81
R1490 vss.t204 vss.t207 1138.81
R1491 vss.t219 vss.t316 1138.81
R1492 vss.t317 vss.t27 1138.81
R1493 vss.t224 vss.t291 1138.81
R1494 vss.t292 vss.t234 1138.81
R1495 vss.t56 vss.t158 1138.81
R1496 vss.t156 vss.t189 1138.81
R1497 vss.t58 vss.t90 1138.81
R1498 vss.t91 vss.t211 1138.81
R1499 vss.t134 vss.t193 1138.81
R1500 vss.t194 vss.t236 1138.81
R1501 vss.t93 vss.t223 1138.81
R1502 vss.t221 vss.t191 1138.81
R1503 vss.t159 vss.t303 1138.81
R1504 vss.t301 vss.t209 1138.81
R1505 vss.t296 vss.t60 1138.81
R1506 vss.t61 vss.t106 1138.81
R1507 vss vss.t355 1134.43
R1508 vss vss.t344 1134.43
R1509 vss vss.t345 1134.43
R1510 vss vss.t354 1134.43
R1511 vss vss.t360 1134.43
R1512 vss vss.t361 1134.43
R1513 vss vss.t11 1134.43
R1514 vss vss.t347 1134.43
R1515 vss vss.t13 1134.43
R1516 vss vss.t12 1134.43
R1517 vss vss.t177 1103.77
R1518 vss vss.t269 1103.77
R1519 vss vss.t169 1103.77
R1520 vss vss.t284 1103.77
R1521 vss vss.t358 1103.77
R1522 vss vss.t244 1103.77
R1523 vss vss.t35 1103.77
R1524 vss vss.t80 1103.77
R1525 vss vss.t149 1103.77
R1526 vss vss.t200 1103.77
R1527 vss.n124 vss.t140 1023.5
R1528 vss.n119 vss.t308 1023.5
R1529 vss.n114 vss.t397 1023.5
R1530 vss.n109 vss.t265 1023.5
R1531 vss.n104 vss.t84 1023.5
R1532 vss.n99 vss.t76 1023.5
R1533 vss.n94 vss.t78 1023.5
R1534 vss.n89 vss.t46 1023.5
R1535 vss.t179 vss.t406 981.133
R1536 vss.t311 vss.t343 981.133
R1537 vss.t267 vss.t39 981.133
R1538 vss.t206 vss.t290 981.133
R1539 vss.t167 vss.t219 981.133
R1540 vss.t316 vss.t370 981.133
R1541 vss.t286 vss.t224 981.133
R1542 vss.t291 vss.t14 981.133
R1543 vss.t356 vss.t56 981.133
R1544 vss.t158 vss.t310 981.133
R1545 vss.t246 vss.t58 981.133
R1546 vss.t90 vss.t44 981.133
R1547 vss.t37 vss.t134 981.133
R1548 vss.t193 vss.t153 981.133
R1549 vss.t82 vss.t93 981.133
R1550 vss.t223 vss.t96 981.133
R1551 vss.t147 vss.t159 981.133
R1552 vss.t303 vss.t175 981.133
R1553 vss.t202 vss.t296 981.133
R1554 vss.t60 vss.t176 981.133
R1555 vss.n83 vss.n2 893.532
R1556 vss.t355 vss.t232 805.931
R1557 vss.n130 vss 805.931
R1558 vss.t344 vss.t5 805.931
R1559 vss vss.n74 805.931
R1560 vss.t345 vss.t321 805.931
R1561 vss vss.n65 805.931
R1562 vss.t354 vss.t271 805.931
R1563 vss vss.n56 805.931
R1564 vss.t360 vss.t215 805.931
R1565 vss vss.n47 805.931
R1566 vss.t361 vss.t127 805.931
R1567 vss vss.n38 805.931
R1568 vss.t11 vss.t198 805.931
R1569 vss vss.n29 805.931
R1570 vss.t347 vss.t399 805.931
R1571 vss vss.n20 805.931
R1572 vss.t13 vss.t29 805.931
R1573 vss vss.n11 805.931
R1574 vss.t12 vss.t329 805.931
R1575 vss vss.n2 805.931
R1576 vss.n7 vss.n5 805.874
R1577 vss.n16 vss.n14 805.874
R1578 vss.n25 vss.n23 805.874
R1579 vss.n34 vss.n32 805.874
R1580 vss.n43 vss.n41 805.874
R1581 vss.n52 vss.n50 805.874
R1582 vss.n61 vss.n59 805.874
R1583 vss.n70 vss.n68 805.874
R1584 vss.n79 vss.n77 805.874
R1585 vss.n84 vss.t145 752.856
R1586 vss.t343 vss.t393 735.85
R1587 vss.t290 vss.t165 735.85
R1588 vss.t370 vss.t154 735.85
R1589 vss.t14 vss.t151 735.85
R1590 vss.t310 vss.t288 735.85
R1591 vss.t44 vss.t171 735.85
R1592 vss.t153 vss.t143 735.85
R1593 vss.t96 vss.t348 735.85
R1594 vss.t175 vss.t33 735.85
R1595 vss.t176 vss.t331 735.85
R1596 vss.t125 vss.t238 593.802
R1597 vss.t262 vss.t323 593.802
R1598 vss.t363 vss.t242 593.802
R1599 vss.t116 vss.t240 593.802
R1600 vss.t279 vss.t408 593.802
R1601 vss.t386 vss.t217 593.802
R1602 vss.t15 vss.t48 593.802
R1603 vss.t378 vss.t325 593.802
R1604 vss.t72 vss.t314 593.802
R1605 vss.n128 vss.n1 533.692
R1606 vss.t232 vss 512.466
R1607 vss.t5 vss 512.466
R1608 vss.t321 vss 512.466
R1609 vss.t271 vss 512.466
R1610 vss.t215 vss 512.466
R1611 vss.t127 vss 512.466
R1612 vss.t198 vss 512.466
R1613 vss.t399 vss 512.466
R1614 vss.t29 vss 512.466
R1615 vss.t329 vss 512.466
R1616 vss.t294 vss 508.087
R1617 vss.t104 vss 508.087
R1618 vss.t140 vss 508.087
R1619 vss.t207 vss 508.087
R1620 vss.t308 vss 508.087
R1621 vss.t27 vss 508.087
R1622 vss.t397 vss 508.087
R1623 vss.t234 vss 508.087
R1624 vss.t265 vss 508.087
R1625 vss.t189 vss 508.087
R1626 vss.t84 vss 508.087
R1627 vss.t211 vss 508.087
R1628 vss.t76 vss 508.087
R1629 vss.t236 vss 508.087
R1630 vss.t78 vss 508.087
R1631 vss.t191 vss 508.087
R1632 vss.t46 vss 508.087
R1633 vss.t209 vss 508.087
R1634 vss.t106 vss 508.087
R1635 vss.t145 vss 491.714
R1636 vss.n130 vss.n129 490.567
R1637 vss.n123 vss.n74 490.567
R1638 vss.n118 vss.n65 490.567
R1639 vss.n113 vss.n56 490.567
R1640 vss.n108 vss.n47 490.567
R1641 vss.n103 vss.n38 490.567
R1642 vss.n98 vss.n29 490.567
R1643 vss.n93 vss.n20 490.567
R1644 vss.n88 vss.n11 490.567
R1645 vss vss.n0 466.558
R1646 vss.n86 vss 408.238
R1647 vss.n91 vss 408.238
R1648 vss.n96 vss 408.238
R1649 vss.n101 vss 408.238
R1650 vss.n106 vss 408.238
R1651 vss.n111 vss 408.238
R1652 vss.n116 vss 408.238
R1653 vss.n121 vss 408.238
R1654 vss.n126 vss 408.238
R1655 vss.n128 vss.t294 376.685
R1656 vss.n303 vss.t0 376.428
R1657 vss.t337 vss.t383 349.918
R1658 vss.t238 vss 307.505
R1659 vss.t323 vss 307.505
R1660 vss.t242 vss 307.505
R1661 vss.t240 vss 307.505
R1662 vss.t408 vss 307.505
R1663 vss.t217 vss 307.505
R1664 vss.t48 vss 307.505
R1665 vss.t325 vss 307.505
R1666 vss.t314 vss 307.505
R1667 vss vss.t337 307.505
R1668 vss.t383 vss 307.505
R1669 vss.n8 vss.n7 265.091
R1670 vss.n17 vss.n16 265.091
R1671 vss.n26 vss.n25 265.091
R1672 vss.n35 vss.n34 265.091
R1673 vss.n44 vss.n43 265.091
R1674 vss.n53 vss.n52 265.091
R1675 vss.n62 vss.n61 265.091
R1676 vss.n71 vss.n70 265.091
R1677 vss.n80 vss.n79 265.091
R1678 vss.n87 vss.t123 245.766
R1679 vss.n92 vss.t258 245.766
R1680 vss.n97 vss.t368 245.766
R1681 vss.n102 vss.t114 245.766
R1682 vss.n107 vss.t281 245.766
R1683 vss.n112 vss.t388 245.766
R1684 vss.n117 vss.t18 245.766
R1685 vss.n122 vss.t376 245.766
R1686 vss.n127 vss.t70 245.766
R1687 vss.n84 vss.n5 233.28
R1688 vss vss.n8 222.675
R1689 vss vss.n17 222.675
R1690 vss vss.n26 222.675
R1691 vss vss.n35 222.675
R1692 vss vss.n44 222.675
R1693 vss vss.n53 222.675
R1694 vss vss.n62 222.675
R1695 vss vss.n71 222.675
R1696 vss vss.n80 222.675
R1697 vss.n303 vss.t404 222.173
R1698 vss.t88 vss.n302 214.308
R1699 vss vss.t249 212.072
R1700 vss vss.t42 212.072
R1701 vss vss.t131 212.072
R1702 vss vss.t298 212.072
R1703 vss vss.t98 212.072
R1704 vss vss.t227 212.072
R1705 vss vss.t109 212.072
R1706 vss vss.t102 212.072
R1707 vss vss.t352 212.072
R1708 vss.n88 vss.t185 176.952
R1709 vss.n93 vss.t23 176.952
R1710 vss.n98 vss.t52 176.952
R1711 vss.n103 vss.t304 176.952
R1712 vss.n108 vss.t255 176.952
R1713 vss.n113 vss.t136 176.952
R1714 vss.n118 vss.t7 176.952
R1715 vss.n123 vss.t161 176.952
R1716 vss.n129 vss.t63 176.952
R1717 vss.t336 vss.t342 157.291
R1718 vss.t339 vss.t335 157.291
R1719 vss.t121 vss.t124 157.291
R1720 vss.t260 vss.t264 157.291
R1721 vss.t367 vss.t369 157.291
R1722 vss.t113 vss.t115 157.291
R1723 vss.t276 vss.t278 157.291
R1724 vss.t391 vss.t385 157.291
R1725 vss.t21 vss.t22 157.291
R1726 vss.t375 vss.t377 157.291
R1727 vss.t68 vss.t71 157.291
R1728 vss.n302 vss.t86 147.459
R1729 vss.t122 vss.t327 133.696
R1730 vss.t261 vss.t31 133.696
R1731 vss.t366 vss.t401 133.696
R1732 vss.t111 vss.t196 133.696
R1733 vss.t277 vss.t129 133.696
R1734 vss.t392 vss.t213 133.696
R1735 vss.t20 vss.t273 133.696
R1736 vss.t373 vss.t319 133.696
R1737 vss.t69 vss.t3 133.696
R1738 vss.t327 vss.n86 131.731
R1739 vss.t31 vss.n91 131.731
R1740 vss.t401 vss.n96 131.731
R1741 vss.t196 vss.n101 131.731
R1742 vss.t129 vss.n106 131.731
R1743 vss.t213 vss.n111 131.731
R1744 vss.t273 vss.n116 131.731
R1745 vss.t319 vss.n121 131.731
R1746 vss.t3 vss.n126 131.731
R1747 vss.t2 vss.t341 129.764
R1748 vss.t341 vss.t333 125.832
R1749 vss.t120 vss.t95 125.832
R1750 vss.t257 vss.t403 125.832
R1751 vss.t365 vss.t75 125.832
R1752 vss.t118 vss.t275 125.832
R1753 vss.t283 vss.t231 125.832
R1754 vss.t390 vss.t142 125.832
R1755 vss.t17 vss.t45 125.832
R1756 vss.t380 vss.t100 125.832
R1757 vss.t74 vss.t350 125.832
R1758 vss.t340 vss.t346 121.9
R1759 vss.t119 vss.t181 121.9
R1760 vss.t259 vss.t371 121.9
R1761 vss.t362 vss.t395 121.9
R1762 vss.t112 vss.t381 121.9
R1763 vss.t282 vss.t229 121.9
R1764 vss.t389 vss.t251 121.9
R1765 vss.t19 vss.t187 121.9
R1766 vss.t374 vss.t50 121.9
R1767 vss.t67 vss.t173 121.9
R1768 vss.n89 vss.n14 111.338
R1769 vss.n94 vss.n23 111.338
R1770 vss.n99 vss.n32 111.338
R1771 vss.n104 vss.n41 111.338
R1772 vss.n109 vss.n50 111.338
R1773 vss.n114 vss.n59 111.338
R1774 vss.n119 vss.n68 111.338
R1775 vss.n124 vss.n77 111.338
R1776 vss.t183 vss.t119 98.3066
R1777 vss.t25 vss.t259 98.3066
R1778 vss.t54 vss.t362 98.3066
R1779 vss.t306 vss.t112 98.3066
R1780 vss.t253 vss.t282 98.3066
R1781 vss.t138 vss.t389 98.3066
R1782 vss.t9 vss.t19 98.3066
R1783 vss.t163 vss.t374 98.3066
R1784 vss.t65 vss.t67 98.3066
R1785 vss.t249 vss.t125 95.4328
R1786 vss.t42 vss.t262 95.4328
R1787 vss.t131 vss.t363 95.4328
R1788 vss.t298 vss.t116 95.4328
R1789 vss.t98 vss.t279 95.4328
R1790 vss.t227 vss.t386 95.4328
R1791 vss.t109 vss.t15 95.4328
R1792 vss.t102 vss.t378 95.4328
R1793 vss.t352 vss.t72 95.4328
R1794 vss.t248 vss.t120 94.3744
R1795 vss.t41 vss.t257 94.3744
R1796 vss.t133 vss.t365 94.3744
R1797 vss.t300 vss.t118 94.3744
R1798 vss.t97 vss.t283 94.3744
R1799 vss.t226 vss.t390 94.3744
R1800 vss.t108 vss.t17 94.3744
R1801 vss.t101 vss.t380 94.3744
R1802 vss.t351 vss.t74 94.3744
R1803 vss.n83 vss.t86 86.5099
R1804 vss.t124 vss.t248 62.9164
R1805 vss.t264 vss.t41 62.9164
R1806 vss.t369 vss.t133 62.9164
R1807 vss.t115 vss.t300 62.9164
R1808 vss.t278 vss.t97 62.9164
R1809 vss.t385 vss.t226 62.9164
R1810 vss.t22 vss.t108 62.9164
R1811 vss.t377 vss.t101 62.9164
R1812 vss.t71 vss.t351 62.9164
R1813 vss.t123 vss.t183 58.9842
R1814 vss.t258 vss.t25 58.9842
R1815 vss.t368 vss.t54 58.9842
R1816 vss.t114 vss.t306 58.9842
R1817 vss.t281 vss.t253 58.9842
R1818 vss.t388 vss.t138 58.9842
R1819 vss.t18 vss.t9 58.9842
R1820 vss.t376 vss.t163 58.9842
R1821 vss.t70 vss.t65 58.9842
R1822 vss.t185 vss.n87 57.018
R1823 vss.t23 vss.n92 57.018
R1824 vss.t52 vss.n97 57.018
R1825 vss.t304 vss.n102 57.018
R1826 vss.t255 vss.n107 57.018
R1827 vss.t136 vss.n112 57.018
R1828 vss.t7 vss.n117 57.018
R1829 vss.t161 vss.n122 57.018
R1830 vss.t63 vss.n127 57.018
R1831 vss.t404 vss.t340 43.2552
R1832 vss.t346 vss.t339 35.3907
R1833 vss.t181 vss.t121 35.3907
R1834 vss.t371 vss.t260 35.3907
R1835 vss.t395 vss.t367 35.3907
R1836 vss.t381 vss.t113 35.3907
R1837 vss.t229 vss.t276 35.3907
R1838 vss.t251 vss.t391 35.3907
R1839 vss.t187 vss.t21 35.3907
R1840 vss.t50 vss.t375 35.3907
R1841 vss.t173 vss.t68 35.3907
R1842 vss.t0 vss 31.8113
R1843 vss.t342 vss.t88 31.4585
R1844 vss.t333 vss.t336 31.4585
R1845 vss.t95 vss.t122 31.4585
R1846 vss.t403 vss.t261 31.4585
R1847 vss.t75 vss.t366 31.4585
R1848 vss.t275 vss.t111 31.4585
R1849 vss.t231 vss.t277 31.4585
R1850 vss.t142 vss.t392 31.4585
R1851 vss.t45 vss.t20 31.4585
R1852 vss.t100 vss.t373 31.4585
R1853 vss.t350 vss.t69 31.4585
R1854 vss.t335 vss.t2 27.5262
R1855 vss.n305 vss.n0 21.2077
R1856 vss.n299 vss.t405 8.79702
R1857 vss.n138 vss.t394 8.79702
R1858 vss.n144 vss.t4 8.79702
R1859 vss.n155 vss.t166 8.79702
R1860 vss.n161 vss.t320 8.79702
R1861 vss.n172 vss.t155 8.79702
R1862 vss.n178 vss.t274 8.79702
R1863 vss.n189 vss.t152 8.79702
R1864 vss.n195 vss.t214 8.79702
R1865 vss.n206 vss.t289 8.79702
R1866 vss.n212 vss.t130 8.79702
R1867 vss.n223 vss.t172 8.79702
R1868 vss.n229 vss.t197 8.79702
R1869 vss.n240 vss.t144 8.79702
R1870 vss.n246 vss.t402 8.79702
R1871 vss.n257 vss.t349 8.79702
R1872 vss.n263 vss.t32 8.79702
R1873 vss.n274 vss.t34 8.79702
R1874 vss.n280 vss.t328 8.79702
R1875 vss.n291 vss.t332 8.79702
R1876 vss.n297 vss.n296 6.40811
R1877 vss.n139 vss.n131 6.40811
R1878 vss.n146 vss.n81 6.40811
R1879 vss.n156 vss.n75 6.40811
R1880 vss.n163 vss.n72 6.40811
R1881 vss.n173 vss.n66 6.40811
R1882 vss.n180 vss.n63 6.40811
R1883 vss.n190 vss.n57 6.40811
R1884 vss.n197 vss.n54 6.40811
R1885 vss.n207 vss.n48 6.40811
R1886 vss.n214 vss.n45 6.40811
R1887 vss.n224 vss.n39 6.40811
R1888 vss.n231 vss.n36 6.40811
R1889 vss.n241 vss.n30 6.40811
R1890 vss.n248 vss.n27 6.40811
R1891 vss.n258 vss.n21 6.40811
R1892 vss.n265 vss.n18 6.40811
R1893 vss.n275 vss.n12 6.40811
R1894 vss.n282 vss.n9 6.40811
R1895 vss.n292 vss.n3 6.40811
R1896 vss.n137 vss.n132 6.4042
R1897 vss.n143 vss.n82 6.4042
R1898 vss.n154 vss.n76 6.4042
R1899 vss.n160 vss.n73 6.4042
R1900 vss.n171 vss.n67 6.4042
R1901 vss.n177 vss.n64 6.4042
R1902 vss.n188 vss.n58 6.4042
R1903 vss.n194 vss.n55 6.4042
R1904 vss.n205 vss.n49 6.4042
R1905 vss.n211 vss.n46 6.4042
R1906 vss.n222 vss.n40 6.4042
R1907 vss.n228 vss.n37 6.4042
R1908 vss.n239 vss.n31 6.4042
R1909 vss.n245 vss.n28 6.4042
R1910 vss.n256 vss.n22 6.4042
R1911 vss.n262 vss.n19 6.4042
R1912 vss.n273 vss.n13 6.4042
R1913 vss.n279 vss.n10 6.4042
R1914 vss.n290 vss.n4 6.4042
R1915 vss.n300 vss.n295 6.4042
R1916 vss.n147 vss.n80 5.28469
R1917 vss.n164 vss.n71 5.28469
R1918 vss.n181 vss.n62 5.28469
R1919 vss.n198 vss.n53 5.28469
R1920 vss.n215 vss.n44 5.28469
R1921 vss.n232 vss.n35 5.28469
R1922 vss.n249 vss.n26 5.28469
R1923 vss.n266 vss.n17 5.28469
R1924 vss.n283 vss.n8 5.28469
R1925 vss.n307 vss.n0 5.28469
R1926 vss.n134 vss.t295 4.63989
R1927 vss.n136 vss.t178 4.63989
R1928 vss.n141 vss.t64 4.63989
R1929 vss.n145 vss.t73 4.63989
R1930 vss.n151 vss.t141 4.63989
R1931 vss.n153 vss.t270 4.63989
R1932 vss.n158 vss.t162 4.63989
R1933 vss.n162 vss.t379 4.63989
R1934 vss.n168 vss.t309 4.63989
R1935 vss.n170 vss.t170 4.63989
R1936 vss.n175 vss.t8 4.63989
R1937 vss.n179 vss.t16 4.63989
R1938 vss.n185 vss.t398 4.63989
R1939 vss.n187 vss.t285 4.63989
R1940 vss.n192 vss.t137 4.63989
R1941 vss.n196 vss.t387 4.63989
R1942 vss.n202 vss.t266 4.63989
R1943 vss.n204 vss.t359 4.63989
R1944 vss.n209 vss.t256 4.63989
R1945 vss.n213 vss.t280 4.63989
R1946 vss.n219 vss.t85 4.63989
R1947 vss.n221 vss.t245 4.63989
R1948 vss.n226 vss.t305 4.63989
R1949 vss.n230 vss.t117 4.63989
R1950 vss.n236 vss.t77 4.63989
R1951 vss.n238 vss.t36 4.63989
R1952 vss.n243 vss.t53 4.63989
R1953 vss.n247 vss.t364 4.63989
R1954 vss.n253 vss.t79 4.63989
R1955 vss.n255 vss.t81 4.63989
R1956 vss.n260 vss.t24 4.63989
R1957 vss.n264 vss.t263 4.63989
R1958 vss.n270 vss.t47 4.63989
R1959 vss.n272 vss.t150 4.63989
R1960 vss.n277 vss.t186 4.63989
R1961 vss.n281 vss.t126 4.63989
R1962 vss.n287 vss.t146 4.63989
R1963 vss.n289 vss.t201 4.63989
R1964 vss.n294 vss.t87 4.63989
R1965 vss.n298 vss.t338 4.63989
R1966 vss.n135 vss.t233 4.51271
R1967 vss.n152 vss.t6 4.51271
R1968 vss.n169 vss.t322 4.51271
R1969 vss.n186 vss.t272 4.51271
R1970 vss.n203 vss.t216 4.51271
R1971 vss.n220 vss.t128 4.51271
R1972 vss.n237 vss.t199 4.51271
R1973 vss.n254 vss.t400 4.51271
R1974 vss.n271 vss.t30 4.51271
R1975 vss.n288 vss.t330 4.51271
R1976 vss.n296 vss.t1 3.9605
R1977 vss.n131 vss.t313 3.9605
R1978 vss.n81 vss.t353 3.9605
R1979 vss.n75 vss.t205 3.9605
R1980 vss.n72 vss.t103 3.9605
R1981 vss.n66 vss.t318 3.9605
R1982 vss.n63 vss.t110 3.9605
R1983 vss.n57 vss.t293 3.9605
R1984 vss.n54 vss.t228 3.9605
R1985 vss.n48 vss.t157 3.9605
R1986 vss.n45 vss.t99 3.9605
R1987 vss.n39 vss.t92 3.9605
R1988 vss.n36 vss.t299 3.9605
R1989 vss.n30 vss.t195 3.9605
R1990 vss.n27 vss.t132 3.9605
R1991 vss.n21 vss.t222 3.9605
R1992 vss.n18 vss.t43 3.9605
R1993 vss.n12 vss.t302 3.9605
R1994 vss.n9 vss.t250 3.9605
R1995 vss.n3 vss.t62 3.9605
R1996 vss.n306 vss.n305 3.6294
R1997 vss.n133 vss.n1 3.6294
R1998 vss.n140 vss.n130 3.6294
R1999 vss.n150 vss.n77 3.6294
R2000 vss.n157 vss.n74 3.6294
R2001 vss.n167 vss.n68 3.6294
R2002 vss.n174 vss.n65 3.6294
R2003 vss.n184 vss.n59 3.6294
R2004 vss.n191 vss.n56 3.6294
R2005 vss.n201 vss.n50 3.6294
R2006 vss.n208 vss.n47 3.6294
R2007 vss.n218 vss.n41 3.6294
R2008 vss.n225 vss.n38 3.6294
R2009 vss.n235 vss.n32 3.6294
R2010 vss.n242 vss.n29 3.6294
R2011 vss.n252 vss.n23 3.6294
R2012 vss.n259 vss.n20 3.6294
R2013 vss.n269 vss.n14 3.6294
R2014 vss.n276 vss.n11 3.6294
R2015 vss.n286 vss.n5 3.6294
R2016 vss.n293 vss.n2 3.6294
R2017 vss.n7 vss.n6 3.46717
R2018 vss.n16 vss.n15 3.46717
R2019 vss.n25 vss.n24 3.46717
R2020 vss.n34 vss.n33 3.46717
R2021 vss.n43 vss.n42 3.46717
R2022 vss.n52 vss.n51 3.46717
R2023 vss.n61 vss.n60 3.46717
R2024 vss.n70 vss.n69 3.46717
R2025 vss.n79 vss.n78 3.46717
R2026 vss.n132 vss.t180 2.07392
R2027 vss.n132 vss.t407 2.07392
R2028 vss.n82 vss.t66 2.07392
R2029 vss.n82 vss.t174 2.07392
R2030 vss.n76 vss.t268 2.07392
R2031 vss.n76 vss.t40 2.07392
R2032 vss.n73 vss.t164 2.07392
R2033 vss.n73 vss.t51 2.07392
R2034 vss.n67 vss.t168 2.07392
R2035 vss.n67 vss.t220 2.07392
R2036 vss.n64 vss.t10 2.07392
R2037 vss.n64 vss.t188 2.07392
R2038 vss.n58 vss.t287 2.07392
R2039 vss.n58 vss.t225 2.07392
R2040 vss.n55 vss.t139 2.07392
R2041 vss.n55 vss.t252 2.07392
R2042 vss.n49 vss.t357 2.07392
R2043 vss.n49 vss.t57 2.07392
R2044 vss.n46 vss.t254 2.07392
R2045 vss.n46 vss.t230 2.07392
R2046 vss.n40 vss.t247 2.07392
R2047 vss.n40 vss.t59 2.07392
R2048 vss.n37 vss.t307 2.07392
R2049 vss.n37 vss.t382 2.07392
R2050 vss.n31 vss.t38 2.07392
R2051 vss.n31 vss.t135 2.07392
R2052 vss.n28 vss.t55 2.07392
R2053 vss.n28 vss.t396 2.07392
R2054 vss.n22 vss.t83 2.07392
R2055 vss.n22 vss.t94 2.07392
R2056 vss.n19 vss.t26 2.07392
R2057 vss.n19 vss.t372 2.07392
R2058 vss.n13 vss.t148 2.07392
R2059 vss.n13 vss.t160 2.07392
R2060 vss.n10 vss.t184 2.07392
R2061 vss.n10 vss.t182 2.07392
R2062 vss.n4 vss.t203 2.07392
R2063 vss.n4 vss.t297 2.07392
R2064 vss.n295 vss.t89 2.07392
R2065 vss.n295 vss.t334 2.07392
R2066 vss.n296 vss.t384 1.84987
R2067 vss.n131 vss.t105 1.84987
R2068 vss.n81 vss.t315 1.84987
R2069 vss.n75 vss.t208 1.84987
R2070 vss.n72 vss.t326 1.84987
R2071 vss.n66 vss.t28 1.84987
R2072 vss.n63 vss.t49 1.84987
R2073 vss.n57 vss.t235 1.84987
R2074 vss.n54 vss.t218 1.84987
R2075 vss.n48 vss.t190 1.84987
R2076 vss.n45 vss.t409 1.84987
R2077 vss.n39 vss.t212 1.84987
R2078 vss.n36 vss.t241 1.84987
R2079 vss.n30 vss.t237 1.84987
R2080 vss.n27 vss.t243 1.84987
R2081 vss.n21 vss.t192 1.84987
R2082 vss.n18 vss.t324 1.84987
R2083 vss.n12 vss.t210 1.84987
R2084 vss.n9 vss.t239 1.84987
R2085 vss.n3 vss.t107 1.84987
R2086 vss.n302 vss 1.48621
R2087 vss.n87 vss 1.48621
R2088 vss.n92 vss 1.48621
R2089 vss.n97 vss 1.48621
R2090 vss.n102 vss 1.48621
R2091 vss.n107 vss 1.48621
R2092 vss.n112 vss 1.48621
R2093 vss.n117 vss 1.48621
R2094 vss.n122 vss 1.48621
R2095 vss.n127 vss 1.48621
R2096 vss.n142 vss 0.7205
R2097 vss.n159 vss 0.7205
R2098 vss.n176 vss 0.7205
R2099 vss.n193 vss 0.7205
R2100 vss.n210 vss 0.7205
R2101 vss.n227 vss 0.7205
R2102 vss.n244 vss 0.7205
R2103 vss.n261 vss 0.7205
R2104 vss.n278 vss 0.7205
R2105 vss vss.n301 0.7205
R2106 vss.n149 vss.n78 0.522085
R2107 vss.n166 vss.n69 0.522085
R2108 vss.n183 vss.n60 0.522085
R2109 vss.n200 vss.n51 0.522085
R2110 vss.n217 vss.n42 0.522085
R2111 vss.n234 vss.n33 0.522085
R2112 vss.n251 vss.n24 0.522085
R2113 vss.n268 vss.n15 0.522085
R2114 vss.n285 vss.n6 0.522085
R2115 vss.n148 vss.n78 0.2471
R2116 vss.n165 vss.n69 0.2471
R2117 vss.n182 vss.n60 0.2471
R2118 vss.n199 vss.n51 0.2471
R2119 vss.n216 vss.n42 0.2471
R2120 vss.n233 vss.n33 0.2471
R2121 vss.n250 vss.n24 0.2471
R2122 vss.n267 vss.n15 0.2471
R2123 vss.n284 vss.n6 0.2471
R2124 vss.n137 vss.n136 0.172371
R2125 vss.n154 vss.n153 0.172371
R2126 vss.n171 vss.n170 0.172371
R2127 vss.n188 vss.n187 0.172371
R2128 vss.n205 vss.n204 0.172371
R2129 vss.n222 vss.n221 0.172371
R2130 vss.n239 vss.n238 0.172371
R2131 vss.n256 vss.n255 0.172371
R2132 vss.n273 vss.n272 0.172371
R2133 vss.n290 vss.n289 0.172371
R2134 vss vss.n137 0.132887
R2135 vss vss.n143 0.132887
R2136 vss vss.n154 0.132887
R2137 vss vss.n160 0.132887
R2138 vss vss.n171 0.132887
R2139 vss vss.n177 0.132887
R2140 vss vss.n188 0.132887
R2141 vss vss.n194 0.132887
R2142 vss vss.n205 0.132887
R2143 vss vss.n211 0.132887
R2144 vss vss.n222 0.132887
R2145 vss vss.n228 0.132887
R2146 vss vss.n239 0.132887
R2147 vss vss.n245 0.132887
R2148 vss vss.n256 0.132887
R2149 vss vss.n262 0.132887
R2150 vss vss.n273 0.132887
R2151 vss vss.n279 0.132887
R2152 vss vss.n290 0.132887
R2153 vss.n300 vss 0.132887
R2154 vss.n143 vss.n142 0.123016
R2155 vss.n160 vss.n159 0.123016
R2156 vss.n177 vss.n176 0.123016
R2157 vss.n194 vss.n193 0.123016
R2158 vss.n211 vss.n210 0.123016
R2159 vss.n228 vss.n227 0.123016
R2160 vss.n245 vss.n244 0.123016
R2161 vss.n262 vss.n261 0.123016
R2162 vss.n279 vss.n278 0.123016
R2163 vss.n138 vss 0.122435
R2164 vss.n155 vss 0.122435
R2165 vss.n172 vss 0.122435
R2166 vss.n189 vss 0.122435
R2167 vss.n206 vss 0.122435
R2168 vss.n223 vss 0.122435
R2169 vss.n240 vss 0.122435
R2170 vss.n257 vss 0.122435
R2171 vss.n274 vss 0.122435
R2172 vss.n291 vss 0.122435
R2173 vss vss.n299 0.122218
R2174 vss.n144 vss 0.121383
R2175 vss.n161 vss 0.121383
R2176 vss.n178 vss 0.121383
R2177 vss.n195 vss 0.121383
R2178 vss.n212 vss 0.121383
R2179 vss.n229 vss 0.121383
R2180 vss.n246 vss 0.121383
R2181 vss.n263 vss 0.121383
R2182 vss.n280 vss 0.121383
R2183 vss vss.n139 0.118952
R2184 vss vss.n156 0.118952
R2185 vss vss.n173 0.118952
R2186 vss vss.n190 0.118952
R2187 vss vss.n207 0.118952
R2188 vss vss.n224 0.118952
R2189 vss vss.n241 0.118952
R2190 vss vss.n258 0.118952
R2191 vss vss.n275 0.118952
R2192 vss vss.n292 0.118952
R2193 vss.n139 vss.n138 0.11779
R2194 vss.n156 vss.n155 0.11779
R2195 vss.n173 vss.n172 0.11779
R2196 vss.n190 vss.n189 0.11779
R2197 vss.n207 vss.n206 0.11779
R2198 vss.n224 vss.n223 0.11779
R2199 vss.n241 vss.n240 0.11779
R2200 vss.n258 vss.n257 0.11779
R2201 vss.n275 vss.n274 0.11779
R2202 vss.n292 vss.n291 0.11779
R2203 vss vss.n134 0.102694
R2204 vss vss.n151 0.102694
R2205 vss vss.n168 0.102694
R2206 vss vss.n185 0.102694
R2207 vss vss.n202 0.102694
R2208 vss vss.n219 0.102694
R2209 vss vss.n236 0.102694
R2210 vss vss.n253 0.102694
R2211 vss vss.n270 0.102694
R2212 vss vss.n287 0.102694
R2213 vss.n301 vss.n300 0.0963064
R2214 vss vss.n133 0.0957258
R2215 vss vss.n150 0.0957258
R2216 vss vss.n167 0.0957258
R2217 vss vss.n184 0.0957258
R2218 vss vss.n201 0.0957258
R2219 vss vss.n218 0.0957258
R2220 vss vss.n235 0.0957258
R2221 vss vss.n252 0.0957258
R2222 vss vss.n269 0.0957258
R2223 vss vss.n286 0.0957258
R2224 vss.n301 vss.n294 0.0765645
R2225 vss.n299 vss.n298 0.06971
R2226 vss.n135 vss 0.0605968
R2227 vss.n152 vss 0.0605968
R2228 vss.n169 vss 0.0605968
R2229 vss.n186 vss 0.0605968
R2230 vss.n203 vss 0.0605968
R2231 vss.n220 vss 0.0605968
R2232 vss.n237 vss 0.0605968
R2233 vss.n254 vss 0.0605968
R2234 vss.n271 vss 0.0605968
R2235 vss.n288 vss 0.0605968
R2236 vss vss.n307 0.05612
R2237 vss.n141 vss.n140 0.0515968
R2238 vss.n158 vss.n157 0.0515968
R2239 vss.n175 vss.n174 0.0515968
R2240 vss.n192 vss.n191 0.0515968
R2241 vss.n209 vss.n208 0.0515968
R2242 vss.n226 vss.n225 0.0515968
R2243 vss.n243 vss.n242 0.0515968
R2244 vss.n260 vss.n259 0.0515968
R2245 vss.n277 vss.n276 0.0515968
R2246 vss.n294 vss.n293 0.0515968
R2247 vss.n142 vss.n141 0.0498548
R2248 vss.n159 vss.n158 0.0498548
R2249 vss.n176 vss.n175 0.0498548
R2250 vss.n193 vss.n192 0.0498548
R2251 vss.n210 vss.n209 0.0498548
R2252 vss.n227 vss.n226 0.0498548
R2253 vss.n244 vss.n243 0.0498548
R2254 vss.n261 vss.n260 0.0498548
R2255 vss.n278 vss.n277 0.0498548
R2256 vss.n134 vss 0.044629
R2257 vss.n151 vss 0.044629
R2258 vss.n168 vss 0.044629
R2259 vss.n185 vss 0.044629
R2260 vss.n202 vss 0.044629
R2261 vss.n219 vss 0.044629
R2262 vss.n236 vss 0.044629
R2263 vss.n253 vss 0.044629
R2264 vss.n270 vss 0.044629
R2265 vss.n287 vss 0.044629
R2266 vss.n145 vss.n144 0.043835
R2267 vss.n162 vss.n161 0.043835
R2268 vss.n179 vss.n178 0.043835
R2269 vss.n196 vss.n195 0.043835
R2270 vss.n213 vss.n212 0.043835
R2271 vss.n230 vss.n229 0.043835
R2272 vss.n247 vss.n246 0.043835
R2273 vss.n264 vss.n263 0.043835
R2274 vss.n281 vss.n280 0.043835
R2275 vss.n306 vss 0.04322
R2276 vss.n136 vss.n135 0.0425968
R2277 vss.n153 vss.n152 0.0425968
R2278 vss.n170 vss.n169 0.0425968
R2279 vss.n187 vss.n186 0.0425968
R2280 vss.n204 vss.n203 0.0425968
R2281 vss.n221 vss.n220 0.0425968
R2282 vss.n238 vss.n237 0.0425968
R2283 vss.n255 vss.n254 0.0425968
R2284 vss.n272 vss.n271 0.0425968
R2285 vss.n289 vss.n288 0.0425968
R2286 vss.n147 vss 0.04082
R2287 vss.n164 vss 0.04082
R2288 vss.n181 vss 0.04082
R2289 vss.n198 vss 0.04082
R2290 vss.n215 vss 0.04082
R2291 vss.n232 vss 0.04082
R2292 vss.n249 vss 0.04082
R2293 vss.n266 vss 0.04082
R2294 vss.n283 vss 0.04082
R2295 vss vss.n149 0.037371
R2296 vss vss.n166 0.037371
R2297 vss vss.n183 0.037371
R2298 vss vss.n200 0.037371
R2299 vss vss.n217 0.037371
R2300 vss vss.n234 0.037371
R2301 vss vss.n251 0.037371
R2302 vss vss.n268 0.037371
R2303 vss vss.n285 0.037371
R2304 vss vss.n145 0.02786
R2305 vss vss.n162 0.02786
R2306 vss vss.n179 0.02786
R2307 vss vss.n196 0.02786
R2308 vss vss.n213 0.02786
R2309 vss vss.n230 0.02786
R2310 vss vss.n247 0.02786
R2311 vss vss.n264 0.02786
R2312 vss vss.n281 0.02786
R2313 vss.n298 vss.n297 0.02426
R2314 vss.n148 vss 0.01616
R2315 vss.n165 vss 0.01616
R2316 vss.n182 vss 0.01616
R2317 vss.n199 vss 0.01616
R2318 vss.n216 vss 0.01616
R2319 vss.n233 vss 0.01616
R2320 vss.n250 vss 0.01616
R2321 vss.n267 vss 0.01616
R2322 vss.n284 vss 0.01616
R2323 vss.n146 vss 0.01346
R2324 vss.n163 vss 0.01346
R2325 vss.n180 vss 0.01346
R2326 vss.n197 vss 0.01346
R2327 vss.n214 vss 0.01346
R2328 vss.n231 vss 0.01346
R2329 vss.n248 vss 0.01346
R2330 vss.n265 vss 0.01346
R2331 vss.n282 vss 0.01346
R2332 vss.n149 vss 0.00787419
R2333 vss.n166 vss 0.00787419
R2334 vss.n183 vss 0.00787419
R2335 vss.n200 vss 0.00787419
R2336 vss.n217 vss 0.00787419
R2337 vss.n234 vss 0.00787419
R2338 vss.n251 vss 0.00787419
R2339 vss.n268 vss 0.00787419
R2340 vss.n285 vss 0.00787419
R2341 vss.n297 vss 0.0041
R2342 vss.n133 vss 0.00282258
R2343 vss.n140 vss 0.00282258
R2344 vss.n150 vss 0.00282258
R2345 vss.n157 vss 0.00282258
R2346 vss.n167 vss 0.00282258
R2347 vss.n174 vss 0.00282258
R2348 vss.n184 vss 0.00282258
R2349 vss.n191 vss 0.00282258
R2350 vss.n201 vss 0.00282258
R2351 vss.n208 vss 0.00282258
R2352 vss.n218 vss 0.00282258
R2353 vss.n225 vss 0.00282258
R2354 vss.n235 vss 0.00282258
R2355 vss.n242 vss 0.00282258
R2356 vss.n252 vss 0.00282258
R2357 vss.n259 vss 0.00282258
R2358 vss.n269 vss 0.00282258
R2359 vss.n276 vss 0.00282258
R2360 vss.n286 vss 0.00282258
R2361 vss.n293 vss 0.00282258
R2362 vss vss.n306 0.00194
R2363 vss vss.n148 0.0014
R2364 vss vss.n165 0.0014
R2365 vss vss.n182 0.0014
R2366 vss vss.n199 0.0014
R2367 vss vss.n216 0.0014
R2368 vss vss.n233 0.0014
R2369 vss vss.n250 0.0014
R2370 vss vss.n267 0.0014
R2371 vss vss.n284 0.0014
R2372 vss vss.n147 0.00122
R2373 vss vss.n164 0.00122
R2374 vss vss.n181 0.00122
R2375 vss vss.n198 0.00122
R2376 vss vss.n215 0.00122
R2377 vss vss.n232 0.00122
R2378 vss vss.n249 0.00122
R2379 vss vss.n266 0.00122
R2380 vss vss.n283 0.00122
R2381 vss vss.n146 0.00104
R2382 vss vss.n163 0.00104
R2383 vss vss.n180 0.00104
R2384 vss vss.n197 0.00104
R2385 vss vss.n214 0.00104
R2386 vss vss.n231 0.00104
R2387 vss vss.n248 0.00104
R2388 vss vss.n265 0.00104
R2389 vss vss.n282 0.00104
R2390 vss.n307 vss 0.00086
R2391 BUS[8].n5 BUS[8].t10 15.5918
R2392 BUS[8].n2 BUS[8].n0 15.3751
R2393 BUS[8].n8 BUS[8].n6 15.2168
R2394 BUS[8].n2 BUS[8].n1 15.0151
R2395 BUS[8].n4 BUS[8].n3 15.0151
R2396 BUS[8].n20 BUS[8].n19 14.8568
R2397 BUS[8].n18 BUS[8].n17 14.8568
R2398 BUS[8].n16 BUS[8].n15 14.8568
R2399 BUS[8].n14 BUS[8].n13 14.8568
R2400 BUS[8].n12 BUS[8].n11 14.8568
R2401 BUS[8].n10 BUS[8].n9 14.8568
R2402 BUS[8].n8 BUS[8].n7 14.8568
R2403 BUS[8].n21 BUS[8] 0.921051
R2404 BUS[8].n5 BUS[8].n4 0.8465
R2405 BUS[8].n19 BUS[8].t13 0.4555
R2406 BUS[8].n19 BUS[8].t17 0.4555
R2407 BUS[8].n17 BUS[8].t12 0.4555
R2408 BUS[8].n17 BUS[8].t11 0.4555
R2409 BUS[8].n15 BUS[8].t9 0.4555
R2410 BUS[8].n15 BUS[8].t14 0.4555
R2411 BUS[8].n13 BUS[8].t1 0.4555
R2412 BUS[8].n13 BUS[8].t20 0.4555
R2413 BUS[8].n11 BUS[8].t21 0.4555
R2414 BUS[8].n11 BUS[8].t18 0.4555
R2415 BUS[8].n9 BUS[8].t22 0.4555
R2416 BUS[8].n9 BUS[8].t16 0.4555
R2417 BUS[8].n7 BUS[8].t19 0.4555
R2418 BUS[8].n7 BUS[8].t15 0.4555
R2419 BUS[8].n6 BUS[8].t8 0.4555
R2420 BUS[8].n6 BUS[8].t0 0.4555
R2421 BUS[8].n0 BUS[8].t2 0.41
R2422 BUS[8].n0 BUS[8].t5 0.41
R2423 BUS[8].n1 BUS[8].t6 0.41
R2424 BUS[8].n1 BUS[8].t7 0.41
R2425 BUS[8].n3 BUS[8].t3 0.41
R2426 BUS[8].n3 BUS[8].t4 0.41
R2427 BUS[8].n4 BUS[8].n2 0.3605
R2428 BUS[8].n10 BUS[8].n8 0.3605
R2429 BUS[8].n12 BUS[8].n10 0.3605
R2430 BUS[8].n14 BUS[8].n12 0.3605
R2431 BUS[8].n16 BUS[8].n14 0.3605
R2432 BUS[8].n18 BUS[8].n16 0.3605
R2433 BUS[8].n20 BUS[8].n18 0.3605
R2434 BUS[8].n21 BUS[8].n5 0.14225
R2435 BUS[8].n21 BUS[8].n20 0.111875
R2436 BUS[8] BUS[8].n21 0.044437
R2437 BUS[1].n5 BUS[1].t22 15.5918
R2438 BUS[1].n2 BUS[1].n0 15.3751
R2439 BUS[1].n8 BUS[1].n6 15.2168
R2440 BUS[1].n2 BUS[1].n1 15.0151
R2441 BUS[1].n4 BUS[1].n3 15.0151
R2442 BUS[1].n20 BUS[1].n19 14.8568
R2443 BUS[1].n18 BUS[1].n17 14.8568
R2444 BUS[1].n16 BUS[1].n15 14.8568
R2445 BUS[1].n14 BUS[1].n13 14.8568
R2446 BUS[1].n12 BUS[1].n11 14.8568
R2447 BUS[1].n10 BUS[1].n9 14.8568
R2448 BUS[1].n8 BUS[1].n7 14.8568
R2449 BUS[1].n21 BUS[1] 0.921051
R2450 BUS[1].n5 BUS[1].n4 0.8465
R2451 BUS[1].n19 BUS[1].t20 0.4555
R2452 BUS[1].n19 BUS[1].t7 0.4555
R2453 BUS[1].n17 BUS[1].t3 0.4555
R2454 BUS[1].n17 BUS[1].t9 0.4555
R2455 BUS[1].n15 BUS[1].t18 0.4555
R2456 BUS[1].n15 BUS[1].t5 0.4555
R2457 BUS[1].n13 BUS[1].t6 0.4555
R2458 BUS[1].n13 BUS[1].t4 0.4555
R2459 BUS[1].n11 BUS[1].t21 0.4555
R2460 BUS[1].n11 BUS[1].t19 0.4555
R2461 BUS[1].n9 BUS[1].t0 0.4555
R2462 BUS[1].n9 BUS[1].t10 0.4555
R2463 BUS[1].n7 BUS[1].t11 0.4555
R2464 BUS[1].n7 BUS[1].t1 0.4555
R2465 BUS[1].n6 BUS[1].t2 0.4555
R2466 BUS[1].n6 BUS[1].t8 0.4555
R2467 BUS[1].n0 BUS[1].t14 0.41
R2468 BUS[1].n0 BUS[1].t15 0.41
R2469 BUS[1].n1 BUS[1].t16 0.41
R2470 BUS[1].n1 BUS[1].t12 0.41
R2471 BUS[1].n3 BUS[1].t17 0.41
R2472 BUS[1].n3 BUS[1].t13 0.41
R2473 BUS[1].n4 BUS[1].n2 0.3605
R2474 BUS[1].n10 BUS[1].n8 0.3605
R2475 BUS[1].n12 BUS[1].n10 0.3605
R2476 BUS[1].n14 BUS[1].n12 0.3605
R2477 BUS[1].n16 BUS[1].n14 0.3605
R2478 BUS[1].n18 BUS[1].n16 0.3605
R2479 BUS[1].n20 BUS[1].n18 0.3605
R2480 BUS[1].n21 BUS[1].n5 0.14225
R2481 BUS[1].n21 BUS[1].n20 0.111875
R2482 BUS[1] BUS[1].n21 0.044437
R2483 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.7994
R2484 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R2485 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2486 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R2487 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R2488 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R2489 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R2490 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R2491 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R2492 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R2493 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R2494 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R2495 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R2496 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R2497 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R2498 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R2499 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R2500 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R2501 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R2502 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R2503 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R2504 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R2505 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R2506 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R2507 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R2508 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R2509 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R2510 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R2511 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R2512 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R2513 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R2514 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R2515 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R2516 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R2517 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R2518 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R2519 BUS[3].n5 BUS[3].t21 15.5918
R2520 BUS[3].n2 BUS[3].n0 15.3751
R2521 BUS[3].n8 BUS[3].n6 15.2168
R2522 BUS[3].n2 BUS[3].n1 15.0151
R2523 BUS[3].n4 BUS[3].n3 15.0151
R2524 BUS[3].n20 BUS[3].n19 14.8568
R2525 BUS[3].n18 BUS[3].n17 14.8568
R2526 BUS[3].n16 BUS[3].n15 14.8568
R2527 BUS[3].n14 BUS[3].n13 14.8568
R2528 BUS[3].n12 BUS[3].n11 14.8568
R2529 BUS[3].n10 BUS[3].n9 14.8568
R2530 BUS[3].n8 BUS[3].n7 14.8568
R2531 BUS[3].n21 BUS[3] 0.921051
R2532 BUS[3].n5 BUS[3].n4 0.8465
R2533 BUS[3].n19 BUS[3].t14 0.4555
R2534 BUS[3].n19 BUS[3].t17 0.4555
R2535 BUS[3].n17 BUS[3].t22 0.4555
R2536 BUS[3].n17 BUS[3].t7 0.4555
R2537 BUS[3].n15 BUS[3].t6 0.4555
R2538 BUS[3].n15 BUS[3].t13 0.4555
R2539 BUS[3].n13 BUS[3].t19 0.4555
R2540 BUS[3].n13 BUS[3].t9 0.4555
R2541 BUS[3].n11 BUS[3].t8 0.4555
R2542 BUS[3].n11 BUS[3].t16 0.4555
R2543 BUS[3].n9 BUS[3].t15 0.4555
R2544 BUS[3].n9 BUS[3].t18 0.4555
R2545 BUS[3].n7 BUS[3].t10 0.4555
R2546 BUS[3].n7 BUS[3].t12 0.4555
R2547 BUS[3].n6 BUS[3].t11 0.4555
R2548 BUS[3].n6 BUS[3].t20 0.4555
R2549 BUS[3].n0 BUS[3].t0 0.41
R2550 BUS[3].n0 BUS[3].t4 0.41
R2551 BUS[3].n1 BUS[3].t3 0.41
R2552 BUS[3].n1 BUS[3].t5 0.41
R2553 BUS[3].n3 BUS[3].t1 0.41
R2554 BUS[3].n3 BUS[3].t2 0.41
R2555 BUS[3].n4 BUS[3].n2 0.3605
R2556 BUS[3].n10 BUS[3].n8 0.3605
R2557 BUS[3].n12 BUS[3].n10 0.3605
R2558 BUS[3].n14 BUS[3].n12 0.3605
R2559 BUS[3].n16 BUS[3].n14 0.3605
R2560 BUS[3].n18 BUS[3].n16 0.3605
R2561 BUS[3].n20 BUS[3].n18 0.3605
R2562 BUS[3].n21 BUS[3].n5 0.14225
R2563 BUS[3].n21 BUS[3].n20 0.111875
R2564 BUS[3] BUS[3].n21 0.044437
R2565 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.7994
R2566 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R2567 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R2568 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R2569 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R2570 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R2571 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R2572 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R2573 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R2574 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R2575 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R2576 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R2577 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R2578 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R2579 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2580 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R2581 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R2582 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R2583 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R2584 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R2585 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R2586 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R2587 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R2588 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R2589 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R2590 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R2591 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R2592 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R2593 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R2594 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R2595 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R2596 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R2597 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R2598 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R2599 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R2600 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R2601 phi_2.n17 phi_2.t19 26.4265
R2602 phi_2.n15 phi_2.t9 26.4265
R2603 phi_2.n13 phi_2.t8 26.4265
R2604 phi_2.n11 phi_2.t16 26.4265
R2605 phi_2.n9 phi_2.t12 26.4265
R2606 phi_2.n7 phi_2.t6 26.4265
R2607 phi_2.n5 phi_2.t0 26.4265
R2608 phi_2.n3 phi_2.t15 26.4265
R2609 phi_2.n1 phi_2.t4 26.4265
R2610 phi_2.n0 phi_2.t18 26.4265
R2611 phi_2.n17 phi_2.t2 11.7657
R2612 phi_2.n15 phi_2.t13 11.7657
R2613 phi_2.n13 phi_2.t10 11.7657
R2614 phi_2.n11 phi_2.t5 11.7657
R2615 phi_2.n9 phi_2.t14 11.7657
R2616 phi_2.n7 phi_2.t7 11.7657
R2617 phi_2.n5 phi_2.t3 11.7657
R2618 phi_2.n3 phi_2.t17 11.7657
R2619 phi_2.n1 phi_2.t11 11.7657
R2620 phi_2.n0 phi_2.t1 11.7657
R2621 phi_2.n18 phi_2 9.23499
R2622 phi_2.n16 phi_2 9.23499
R2623 phi_2.n14 phi_2 9.23499
R2624 phi_2.n12 phi_2 9.23499
R2625 phi_2.n10 phi_2 9.23499
R2626 phi_2.n8 phi_2 9.23499
R2627 phi_2.n6 phi_2 9.23499
R2628 phi_2.n4 phi_2 9.23499
R2629 phi_2.n2 phi_2 9.23499
R2630 phi_2 phi_2.n17 8.04257
R2631 phi_2 phi_2.n15 8.04257
R2632 phi_2 phi_2.n13 8.04257
R2633 phi_2 phi_2.n11 8.04257
R2634 phi_2 phi_2.n9 8.04257
R2635 phi_2 phi_2.n7 8.04257
R2636 phi_2 phi_2.n5 8.04257
R2637 phi_2 phi_2.n3 8.04257
R2638 phi_2 phi_2.n1 8.04257
R2639 phi_2 phi_2.n0 8.04257
R2640 phi_2.n2 phi_2 3.0407
R2641 phi_2.n4 phi_2 3.0407
R2642 phi_2.n6 phi_2 3.0407
R2643 phi_2.n8 phi_2 3.0407
R2644 phi_2.n10 phi_2 3.0407
R2645 phi_2.n12 phi_2 3.0407
R2646 phi_2.n14 phi_2 3.0407
R2647 phi_2.n16 phi_2 3.0407
R2648 phi_2.n18 phi_2 3.0407
R2649 phi_2 phi_2.n2 2.5763
R2650 phi_2 phi_2.n4 2.5763
R2651 phi_2 phi_2.n6 2.5763
R2652 phi_2 phi_2.n8 2.5763
R2653 phi_2 phi_2.n10 2.5763
R2654 phi_2 phi_2.n12 2.5763
R2655 phi_2 phi_2.n14 2.5763
R2656 phi_2 phi_2.n16 2.5763
R2657 phi_2 phi_2.n18 2.5763
R2658 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.7994
R2659 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R2660 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R2661 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R2662 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R2663 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R2664 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R2665 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R2666 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R2667 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R2668 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2669 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R2670 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R2671 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R2672 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R2673 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R2674 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R2675 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R2676 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R2677 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R2678 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R2679 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R2680 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R2681 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R2682 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R2683 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R2684 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R2685 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R2686 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R2687 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R2688 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R2689 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R2690 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R2691 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R2692 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R2693 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R2694 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.7994
R2695 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R2696 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R2697 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R2698 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2699 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R2700 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R2701 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R2702 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R2703 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R2704 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R2705 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R2706 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R2707 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R2708 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R2709 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R2710 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R2711 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R2712 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R2713 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R2714 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R2715 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R2716 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R2717 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R2718 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R2719 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R2720 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R2721 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R2722 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R2723 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R2724 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R2725 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R2726 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R2727 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R2728 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R2729 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R2730 BUS[6].n5 BUS[6].t8 15.5918
R2731 BUS[6].n2 BUS[6].n0 15.3751
R2732 BUS[6].n8 BUS[6].n6 15.2168
R2733 BUS[6].n2 BUS[6].n1 15.0151
R2734 BUS[6].n4 BUS[6].n3 15.0151
R2735 BUS[6].n20 BUS[6].n19 14.8568
R2736 BUS[6].n18 BUS[6].n17 14.8568
R2737 BUS[6].n16 BUS[6].n15 14.8568
R2738 BUS[6].n14 BUS[6].n13 14.8568
R2739 BUS[6].n12 BUS[6].n11 14.8568
R2740 BUS[6].n10 BUS[6].n9 14.8568
R2741 BUS[6].n8 BUS[6].n7 14.8568
R2742 BUS[6].n21 BUS[6] 0.921051
R2743 BUS[6].n5 BUS[6].n4 0.8465
R2744 BUS[6].n19 BUS[6].t14 0.4555
R2745 BUS[6].n19 BUS[6].t0 0.4555
R2746 BUS[6].n17 BUS[6].t4 0.4555
R2747 BUS[6].n17 BUS[6].t11 0.4555
R2748 BUS[6].n15 BUS[6].t10 0.4555
R2749 BUS[6].n15 BUS[6].t2 0.4555
R2750 BUS[6].n13 BUS[6].t1 0.4555
R2751 BUS[6].n13 BUS[6].t9 0.4555
R2752 BUS[6].n11 BUS[6].t13 0.4555
R2753 BUS[6].n11 BUS[6].t15 0.4555
R2754 BUS[6].n9 BUS[6].t3 0.4555
R2755 BUS[6].n9 BUS[6].t6 0.4555
R2756 BUS[6].n7 BUS[6].t5 0.4555
R2757 BUS[6].n7 BUS[6].t12 0.4555
R2758 BUS[6].n6 BUS[6].t16 0.4555
R2759 BUS[6].n6 BUS[6].t7 0.4555
R2760 BUS[6].n0 BUS[6].t22 0.41
R2761 BUS[6].n0 BUS[6].t18 0.41
R2762 BUS[6].n1 BUS[6].t17 0.41
R2763 BUS[6].n1 BUS[6].t19 0.41
R2764 BUS[6].n3 BUS[6].t20 0.41
R2765 BUS[6].n3 BUS[6].t21 0.41
R2766 BUS[6].n4 BUS[6].n2 0.3605
R2767 BUS[6].n10 BUS[6].n8 0.3605
R2768 BUS[6].n12 BUS[6].n10 0.3605
R2769 BUS[6].n14 BUS[6].n12 0.3605
R2770 BUS[6].n16 BUS[6].n14 0.3605
R2771 BUS[6].n18 BUS[6].n16 0.3605
R2772 BUS[6].n20 BUS[6].n18 0.3605
R2773 BUS[6].n21 BUS[6].n5 0.14225
R2774 BUS[6].n21 BUS[6].n20 0.111875
R2775 BUS[6] BUS[6].n21 0.044437
R2776 BUS[10].n5 BUS[10].t7 15.5918
R2777 BUS[10].n2 BUS[10].n0 15.3751
R2778 BUS[10].n8 BUS[10].n6 15.2168
R2779 BUS[10].n2 BUS[10].n1 15.0151
R2780 BUS[10].n4 BUS[10].n3 15.0151
R2781 BUS[10].n20 BUS[10].n19 14.8568
R2782 BUS[10].n18 BUS[10].n17 14.8568
R2783 BUS[10].n16 BUS[10].n15 14.8568
R2784 BUS[10].n14 BUS[10].n13 14.8568
R2785 BUS[10].n12 BUS[10].n11 14.8568
R2786 BUS[10].n10 BUS[10].n9 14.8568
R2787 BUS[10].n8 BUS[10].n7 14.8568
R2788 BUS[10].n21 BUS[10] 0.921051
R2789 BUS[10].n5 BUS[10].n4 0.8465
R2790 BUS[10].n19 BUS[10].t12 0.4555
R2791 BUS[10].n19 BUS[10].t20 0.4555
R2792 BUS[10].n17 BUS[10].t16 0.4555
R2793 BUS[10].n17 BUS[10].t15 0.4555
R2794 BUS[10].n15 BUS[10].t8 0.4555
R2795 BUS[10].n15 BUS[10].t21 0.4555
R2796 BUS[10].n13 BUS[10].t10 0.4555
R2797 BUS[10].n13 BUS[10].t6 0.4555
R2798 BUS[10].n11 BUS[10].t22 0.4555
R2799 BUS[10].n11 BUS[10].t13 0.4555
R2800 BUS[10].n9 BUS[10].t14 0.4555
R2801 BUS[10].n9 BUS[10].t17 0.4555
R2802 BUS[10].n7 BUS[10].t18 0.4555
R2803 BUS[10].n7 BUS[10].t19 0.4555
R2804 BUS[10].n6 BUS[10].t9 0.4555
R2805 BUS[10].n6 BUS[10].t11 0.4555
R2806 BUS[10].n0 BUS[10].t5 0.41
R2807 BUS[10].n0 BUS[10].t2 0.41
R2808 BUS[10].n1 BUS[10].t1 0.41
R2809 BUS[10].n1 BUS[10].t4 0.41
R2810 BUS[10].n3 BUS[10].t3 0.41
R2811 BUS[10].n3 BUS[10].t0 0.41
R2812 BUS[10].n4 BUS[10].n2 0.3605
R2813 BUS[10].n10 BUS[10].n8 0.3605
R2814 BUS[10].n12 BUS[10].n10 0.3605
R2815 BUS[10].n14 BUS[10].n12 0.3605
R2816 BUS[10].n16 BUS[10].n14 0.3605
R2817 BUS[10].n18 BUS[10].n16 0.3605
R2818 BUS[10].n20 BUS[10].n18 0.3605
R2819 BUS[10].n21 BUS[10].n5 0.14225
R2820 BUS[10].n21 BUS[10].n20 0.111875
R2821 BUS[10] BUS[10].n21 0.044437
R2822 enable.n18 enable.t10 19.9538
R2823 enable.n16 enable.t11 19.9538
R2824 enable.n14 enable.t4 19.9538
R2825 enable.n12 enable.t8 19.9538
R2826 enable.n10 enable.t17 19.9538
R2827 enable.n8 enable.t19 19.9538
R2828 enable.n6 enable.t5 19.9538
R2829 enable.n4 enable.t15 19.9538
R2830 enable.n2 enable.t0 19.9538
R2831 enable.n0 enable.t7 19.9538
R2832 enable.n18 enable.t2 17.3015
R2833 enable.n16 enable.t3 17.3015
R2834 enable.n14 enable.t14 17.3015
R2835 enable.n12 enable.t18 17.3015
R2836 enable.n10 enable.t6 17.3015
R2837 enable.n8 enable.t12 17.3015
R2838 enable.n6 enable.t16 17.3015
R2839 enable.n4 enable.t9 17.3015
R2840 enable.n2 enable.t13 17.3015
R2841 enable.n0 enable.t1 17.3015
R2842 enable enable.n19 10.8498
R2843 enable.n19 enable.n18 8.0005
R2844 enable.n17 enable.n16 8.0005
R2845 enable.n15 enable.n14 8.0005
R2846 enable.n13 enable.n12 8.0005
R2847 enable.n11 enable.n10 8.0005
R2848 enable.n9 enable.n8 8.0005
R2849 enable.n7 enable.n6 8.0005
R2850 enable.n5 enable.n4 8.0005
R2851 enable.n3 enable.n2 8.0005
R2852 enable.n1 enable.n0 8.0005
R2853 enable enable.n20 6.01421
R2854 enable enable.n21 6.01421
R2855 enable enable.n22 6.01421
R2856 enable enable.n23 6.01421
R2857 enable enable.n24 6.01421
R2858 enable enable.n25 6.01421
R2859 enable enable.n26 6.01421
R2860 enable enable.n27 6.01421
R2861 enable enable.n28 6.01421
R2862 enable.n20 enable.n17 4.8361
R2863 enable.n21 enable.n15 4.8361
R2864 enable.n22 enable.n13 4.8361
R2865 enable.n23 enable.n11 4.8361
R2866 enable.n24 enable.n9 4.8361
R2867 enable.n25 enable.n7 4.8361
R2868 enable.n26 enable.n5 4.8361
R2869 enable.n27 enable.n3 4.8361
R2870 enable.n28 enable.n1 4.8361
R2871 enable.n20 enable 1.07965
R2872 enable.n21 enable 1.07965
R2873 enable.n22 enable 1.07965
R2874 enable.n23 enable 1.07965
R2875 enable.n24 enable 1.07965
R2876 enable.n25 enable 1.07965
R2877 enable.n26 enable 1.07965
R2878 enable.n27 enable 1.07965
R2879 enable.n28 enable 1.07965
R2880 enable.n19 enable 0.00742308
R2881 enable.n17 enable 0.00742308
R2882 enable.n15 enable 0.00742308
R2883 enable.n13 enable 0.00742308
R2884 enable.n11 enable 0.00742308
R2885 enable.n9 enable 0.00742308
R2886 enable.n7 enable 0.00742308
R2887 enable.n5 enable 0.00742308
R2888 enable.n3 enable 0.00742308
R2889 enable.n1 enable 0.00742308
R2890 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.7994
R2891 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R2892 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R2893 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R2894 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R2895 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R2896 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R2897 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R2898 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R2899 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R2900 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R2901 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R2902 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R2903 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R2904 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R2905 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R2906 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R2907 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R2908 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R2909 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R2910 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R2911 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R2912 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R2913 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R2914 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R2915 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R2916 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R2917 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R2918 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R2919 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R2920 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R2921 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R2922 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R2923 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R2924 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R2925 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R2926 BUS[2].n5 BUS[2].t12 15.5918
R2927 BUS[2].n2 BUS[2].n0 15.3751
R2928 BUS[2].n8 BUS[2].n6 15.2168
R2929 BUS[2].n2 BUS[2].n1 15.0151
R2930 BUS[2].n4 BUS[2].n3 15.0151
R2931 BUS[2].n20 BUS[2].n19 14.8568
R2932 BUS[2].n18 BUS[2].n17 14.8568
R2933 BUS[2].n16 BUS[2].n15 14.8568
R2934 BUS[2].n14 BUS[2].n13 14.8568
R2935 BUS[2].n12 BUS[2].n11 14.8568
R2936 BUS[2].n10 BUS[2].n9 14.8568
R2937 BUS[2].n8 BUS[2].n7 14.8568
R2938 BUS[2].n21 BUS[2] 0.921051
R2939 BUS[2].n5 BUS[2].n4 0.8465
R2940 BUS[2].n19 BUS[2].t5 0.4555
R2941 BUS[2].n19 BUS[2].t9 0.4555
R2942 BUS[2].n17 BUS[2].t14 0.4555
R2943 BUS[2].n17 BUS[2].t2 0.4555
R2944 BUS[2].n15 BUS[2].t1 0.4555
R2945 BUS[2].n15 BUS[2].t4 0.4555
R2946 BUS[2].n13 BUS[2].t10 0.4555
R2947 BUS[2].n13 BUS[2].t13 0.4555
R2948 BUS[2].n11 BUS[2].t0 0.4555
R2949 BUS[2].n11 BUS[2].t7 0.4555
R2950 BUS[2].n9 BUS[2].t6 0.4555
R2951 BUS[2].n9 BUS[2].t16 0.4555
R2952 BUS[2].n7 BUS[2].t15 0.4555
R2953 BUS[2].n7 BUS[2].t3 0.4555
R2954 BUS[2].n6 BUS[2].t8 0.4555
R2955 BUS[2].n6 BUS[2].t11 0.4555
R2956 BUS[2].n0 BUS[2].t18 0.41
R2957 BUS[2].n0 BUS[2].t20 0.41
R2958 BUS[2].n1 BUS[2].t19 0.41
R2959 BUS[2].n1 BUS[2].t22 0.41
R2960 BUS[2].n3 BUS[2].t21 0.41
R2961 BUS[2].n3 BUS[2].t17 0.41
R2962 BUS[2].n4 BUS[2].n2 0.3605
R2963 BUS[2].n10 BUS[2].n8 0.3605
R2964 BUS[2].n12 BUS[2].n10 0.3605
R2965 BUS[2].n14 BUS[2].n12 0.3605
R2966 BUS[2].n16 BUS[2].n14 0.3605
R2967 BUS[2].n18 BUS[2].n16 0.3605
R2968 BUS[2].n20 BUS[2].n18 0.3605
R2969 BUS[2].n21 BUS[2].n5 0.14225
R2970 BUS[2].n21 BUS[2].n20 0.111875
R2971 BUS[2] BUS[2].n21 0.044437
R2972 phi_1.n17 phi_1.t2 26.4265
R2973 phi_1.n15 phi_1.t9 26.4265
R2974 phi_1.n13 phi_1.t1 26.4265
R2975 phi_1.n11 phi_1.t12 26.4265
R2976 phi_1.n9 phi_1.t11 26.4265
R2977 phi_1.n7 phi_1.t19 26.4265
R2978 phi_1.n5 phi_1.t16 26.4265
R2979 phi_1.n3 phi_1.t8 26.4265
R2980 phi_1.n1 phi_1.t4 26.4265
R2981 phi_1.n0 phi_1.t18 26.4265
R2982 phi_1.n17 phi_1.t3 11.7657
R2983 phi_1.n15 phi_1.t13 11.7657
R2984 phi_1.n13 phi_1.t5 11.7657
R2985 phi_1.n11 phi_1.t15 11.7657
R2986 phi_1.n9 phi_1.t14 11.7657
R2987 phi_1.n7 phi_1.t7 11.7657
R2988 phi_1.n5 phi_1.t17 11.7657
R2989 phi_1.n3 phi_1.t10 11.7657
R2990 phi_1.n1 phi_1.t6 11.7657
R2991 phi_1.n0 phi_1.t0 11.7657
R2992 phi_1.n18 phi_1 9.56151
R2993 phi_1.n16 phi_1 9.56151
R2994 phi_1.n14 phi_1 9.56151
R2995 phi_1.n12 phi_1 9.56151
R2996 phi_1.n10 phi_1 9.56151
R2997 phi_1.n8 phi_1 9.56151
R2998 phi_1.n6 phi_1 9.56151
R2999 phi_1.n4 phi_1 9.56151
R3000 phi_1.n2 phi_1 9.56151
R3001 phi_1 phi_1.n17 8.04713
R3002 phi_1 phi_1.n15 8.04713
R3003 phi_1 phi_1.n13 8.04713
R3004 phi_1 phi_1.n11 8.04713
R3005 phi_1 phi_1.n9 8.04713
R3006 phi_1 phi_1.n7 8.04713
R3007 phi_1 phi_1.n5 8.04713
R3008 phi_1 phi_1.n3 8.04713
R3009 phi_1 phi_1.n1 8.04713
R3010 phi_1 phi_1.n0 8.04713
R3011 phi_1.n2 phi_1 5.2583
R3012 phi_1.n4 phi_1 5.2583
R3013 phi_1.n6 phi_1 5.2583
R3014 phi_1.n8 phi_1 5.2583
R3015 phi_1.n10 phi_1 5.2583
R3016 phi_1.n12 phi_1 5.2583
R3017 phi_1.n14 phi_1 5.2583
R3018 phi_1.n16 phi_1 5.2583
R3019 phi_1.n18 phi_1 5.2583
R3020 phi_1 phi_1.n2 0.3587
R3021 phi_1 phi_1.n4 0.3587
R3022 phi_1 phi_1.n6 0.3587
R3023 phi_1 phi_1.n8 0.3587
R3024 phi_1 phi_1.n10 0.3587
R3025 phi_1 phi_1.n12 0.3587
R3026 phi_1 phi_1.n14 0.3587
R3027 phi_1 phi_1.n16 0.3587
R3028 phi_1 phi_1.n18 0.3587
R3029 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.7994
R3030 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R3031 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R3032 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R3033 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R3034 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R3035 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R3036 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R3037 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R3038 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R3039 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R3040 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R3041 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R3042 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R3043 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R3044 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R3045 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R3046 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R3047 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R3048 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R3049 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R3050 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R3051 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R3052 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R3053 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R3054 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R3055 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R3056 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R3057 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R3058 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R3059 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R3060 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R3061 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R3062 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R3063 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R3064 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R3065 BUS[4].n5 BUS[4].t15 15.5918
R3066 BUS[4].n2 BUS[4].n0 15.3751
R3067 BUS[4].n8 BUS[4].n6 15.2168
R3068 BUS[4].n2 BUS[4].n1 15.0151
R3069 BUS[4].n4 BUS[4].n3 15.0151
R3070 BUS[4].n20 BUS[4].n19 14.8568
R3071 BUS[4].n18 BUS[4].n17 14.8568
R3072 BUS[4].n16 BUS[4].n15 14.8568
R3073 BUS[4].n14 BUS[4].n13 14.8568
R3074 BUS[4].n12 BUS[4].n11 14.8568
R3075 BUS[4].n10 BUS[4].n9 14.8568
R3076 BUS[4].n8 BUS[4].n7 14.8568
R3077 BUS[4].n21 BUS[4] 0.921051
R3078 BUS[4].n5 BUS[4].n4 0.8465
R3079 BUS[4].n19 BUS[4].t0 0.4555
R3080 BUS[4].n19 BUS[4].t8 0.4555
R3081 BUS[4].n17 BUS[4].t7 0.4555
R3082 BUS[4].n17 BUS[4].t14 0.4555
R3083 BUS[4].n15 BUS[4].t2 0.4555
R3084 BUS[4].n15 BUS[4].t5 0.4555
R3085 BUS[4].n13 BUS[4].t10 0.4555
R3086 BUS[4].n13 BUS[4].t12 0.4555
R3087 BUS[4].n11 BUS[4].t16 0.4555
R3088 BUS[4].n11 BUS[4].t1 0.4555
R3089 BUS[4].n9 BUS[4].t6 0.4555
R3090 BUS[4].n9 BUS[4].t9 0.4555
R3091 BUS[4].n7 BUS[4].t13 0.4555
R3092 BUS[4].n7 BUS[4].t4 0.4555
R3093 BUS[4].n6 BUS[4].t3 0.4555
R3094 BUS[4].n6 BUS[4].t11 0.4555
R3095 BUS[4].n0 BUS[4].t18 0.41
R3096 BUS[4].n0 BUS[4].t19 0.41
R3097 BUS[4].n1 BUS[4].t20 0.41
R3098 BUS[4].n1 BUS[4].t22 0.41
R3099 BUS[4].n3 BUS[4].t21 0.41
R3100 BUS[4].n3 BUS[4].t17 0.41
R3101 BUS[4].n4 BUS[4].n2 0.3605
R3102 BUS[4].n10 BUS[4].n8 0.3605
R3103 BUS[4].n12 BUS[4].n10 0.3605
R3104 BUS[4].n14 BUS[4].n12 0.3605
R3105 BUS[4].n16 BUS[4].n14 0.3605
R3106 BUS[4].n18 BUS[4].n16 0.3605
R3107 BUS[4].n20 BUS[4].n18 0.3605
R3108 BUS[4].n21 BUS[4].n5 0.14225
R3109 BUS[4].n21 BUS[4].n20 0.111875
R3110 BUS[4] BUS[4].n21 0.044437
R3111 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.7994
R3112 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R3113 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R3114 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R3115 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R3116 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R3117 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R3118 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R3119 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R3120 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R3121 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R3122 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R3123 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R3124 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R3125 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R3126 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R3127 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R3128 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R3129 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R3130 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R3131 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R3132 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R3133 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R3134 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R3135 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R3136 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R3137 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R3138 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R3139 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R3140 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R3141 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R3142 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R3143 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R3144 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R3145 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R3146 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R3147 BUS[9].n5 BUS[9].t7 15.5918
R3148 BUS[9].n2 BUS[9].n0 15.3751
R3149 BUS[9].n8 BUS[9].n6 15.2168
R3150 BUS[9].n2 BUS[9].n1 15.0151
R3151 BUS[9].n4 BUS[9].n3 15.0151
R3152 BUS[9].n20 BUS[9].n19 14.8568
R3153 BUS[9].n18 BUS[9].n17 14.8568
R3154 BUS[9].n16 BUS[9].n15 14.8568
R3155 BUS[9].n14 BUS[9].n13 14.8568
R3156 BUS[9].n12 BUS[9].n11 14.8568
R3157 BUS[9].n10 BUS[9].n9 14.8568
R3158 BUS[9].n8 BUS[9].n7 14.8568
R3159 BUS[9].n21 BUS[9] 0.921051
R3160 BUS[9].n5 BUS[9].n4 0.8465
R3161 BUS[9].n19 BUS[9].t13 0.4555
R3162 BUS[9].n19 BUS[9].t15 0.4555
R3163 BUS[9].n17 BUS[9].t5 0.4555
R3164 BUS[9].n17 BUS[9].t2 0.4555
R3165 BUS[9].n15 BUS[9].t9 0.4555
R3166 BUS[9].n15 BUS[9].t1 0.4555
R3167 BUS[9].n13 BUS[9].t14 0.4555
R3168 BUS[9].n13 BUS[9].t22 0.4555
R3169 BUS[9].n11 BUS[9].t6 0.4555
R3170 BUS[9].n11 BUS[9].t10 0.4555
R3171 BUS[9].n9 BUS[9].t3 0.4555
R3172 BUS[9].n9 BUS[9].t8 0.4555
R3173 BUS[9].n7 BUS[9].t4 0.4555
R3174 BUS[9].n7 BUS[9].t11 0.4555
R3175 BUS[9].n6 BUS[9].t12 0.4555
R3176 BUS[9].n6 BUS[9].t0 0.4555
R3177 BUS[9].n0 BUS[9].t21 0.41
R3178 BUS[9].n0 BUS[9].t16 0.41
R3179 BUS[9].n1 BUS[9].t18 0.41
R3180 BUS[9].n1 BUS[9].t20 0.41
R3181 BUS[9].n3 BUS[9].t19 0.41
R3182 BUS[9].n3 BUS[9].t17 0.41
R3183 BUS[9].n4 BUS[9].n2 0.3605
R3184 BUS[9].n10 BUS[9].n8 0.3605
R3185 BUS[9].n12 BUS[9].n10 0.3605
R3186 BUS[9].n14 BUS[9].n12 0.3605
R3187 BUS[9].n16 BUS[9].n14 0.3605
R3188 BUS[9].n18 BUS[9].n16 0.3605
R3189 BUS[9].n20 BUS[9].n18 0.3605
R3190 BUS[9].n21 BUS[9].n5 0.14225
R3191 BUS[9].n21 BUS[9].n20 0.111875
R3192 BUS[9] BUS[9].n21 0.044437
R3193 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.7994
R3194 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R3195 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R3196 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R3197 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R3198 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R3199 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R3200 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R3201 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R3202 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R3203 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R3204 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R3205 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R3206 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R3207 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R3208 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R3209 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R3210 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R3211 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R3212 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R3213 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R3214 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R3215 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R3216 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R3217 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R3218 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R3219 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R3220 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R3221 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R3222 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R3223 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R3224 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R3225 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R3226 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R3227 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R3228 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R3229 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.7994
R3230 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R3231 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.6148
R3232 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R3233 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R3234 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R3235 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R3236 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R3237 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R3238 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R3239 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R3240 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R3241 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R3242 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R3243 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R3244 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R3245 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R3246 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 11.7121
R3247 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 4.63372
R3248 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 3.85252
R3249 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 0.402556
R3250 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R3251 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R3252 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R3253 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R3254 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R3255 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R3256 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R3257 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R3258 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R3259 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R3260 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R3261 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R3262 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R3263 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R3264 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R3265 BUS[7].n5 BUS[7].t6 15.5918
R3266 BUS[7].n2 BUS[7].n0 15.3751
R3267 BUS[7].n8 BUS[7].n6 15.2168
R3268 BUS[7].n2 BUS[7].n1 15.0151
R3269 BUS[7].n4 BUS[7].n3 15.0151
R3270 BUS[7].n20 BUS[7].n19 14.8568
R3271 BUS[7].n18 BUS[7].n17 14.8568
R3272 BUS[7].n16 BUS[7].n15 14.8568
R3273 BUS[7].n14 BUS[7].n13 14.8568
R3274 BUS[7].n12 BUS[7].n11 14.8568
R3275 BUS[7].n10 BUS[7].n9 14.8568
R3276 BUS[7].n8 BUS[7].n7 14.8568
R3277 BUS[7].n21 BUS[7] 0.921051
R3278 BUS[7].n5 BUS[7].n4 0.8465
R3279 BUS[7].n19 BUS[7].t12 0.4555
R3280 BUS[7].n19 BUS[7].t1 0.4555
R3281 BUS[7].n17 BUS[7].t0 0.4555
R3282 BUS[7].n17 BUS[7].t9 0.4555
R3283 BUS[7].n15 BUS[7].t8 0.4555
R3284 BUS[7].n15 BUS[7].t11 0.4555
R3285 BUS[7].n13 BUS[7].t3 0.4555
R3286 BUS[7].n13 BUS[7].t5 0.4555
R3287 BUS[7].n11 BUS[7].t4 0.4555
R3288 BUS[7].n11 BUS[7].t14 0.4555
R3289 BUS[7].n9 BUS[7].t13 0.4555
R3290 BUS[7].n9 BUS[7].t2 0.4555
R3291 BUS[7].n7 BUS[7].t7 0.4555
R3292 BUS[7].n7 BUS[7].t10 0.4555
R3293 BUS[7].n6 BUS[7].t15 0.4555
R3294 BUS[7].n6 BUS[7].t16 0.4555
R3295 BUS[7].n0 BUS[7].t20 0.41
R3296 BUS[7].n0 BUS[7].t22 0.41
R3297 BUS[7].n1 BUS[7].t21 0.41
R3298 BUS[7].n1 BUS[7].t17 0.41
R3299 BUS[7].n3 BUS[7].t18 0.41
R3300 BUS[7].n3 BUS[7].t19 0.41
R3301 BUS[7].n4 BUS[7].n2 0.3605
R3302 BUS[7].n10 BUS[7].n8 0.3605
R3303 BUS[7].n12 BUS[7].n10 0.3605
R3304 BUS[7].n14 BUS[7].n12 0.3605
R3305 BUS[7].n16 BUS[7].n14 0.3605
R3306 BUS[7].n18 BUS[7].n16 0.3605
R3307 BUS[7].n20 BUS[7].n18 0.3605
R3308 BUS[7].n21 BUS[7].n5 0.14225
R3309 BUS[7].n21 BUS[7].n20 0.111875
R3310 BUS[7] BUS[7].n21 0.044437
R3311 d_out.n0 d_out.t2 21.1948
R3312 d_out.n0 d_out.t3 16.0605
R3313 d_out d_out.n3 9.16609
R3314 d_out.n2 d_out.n1 9.0005
R3315 d_out.n1 d_out.n0 8.12012
R3316 d_out.n2 d_out 5.47636
R3317 d_out.n3 d_out.t0 4.5901
R3318 d_out d_out.t1 3.91488
R3319 d_out.n3 d_out 0.150731
R3320 d_out d_out.n2 0.13775
R3321 d_out.n1 d_out 0.00840541
R3322 D_in.n0 D_in.t0 29.4195
R3323 D_in.n0 D_in.t1 11.4372
R3324 D_in D_in.n1 9.95
R3325 D_in.n1 D_in.n0 8.0005
R3326 D_in.n1 D_in 0.102506
C0 a_53720_2002# d_out 0
C1 a_32536_2002# BUS[6] 0.01182f
C2 swmatrix_Tgate_2.gated_control a_59468_1577# 0
C3 a_47480_2002# a_47380_1577# 0
C4 swmatrix_Tgate_6.gated_control phi_1 0.01084f
C5 a_46620_1580# a_46988_1577# 0.00194f
C6 a_43688_1562# BUS[8] 0.00406f
C7 a_27900_1580# swmatrix_Tgate_5.gated_control 0.00668f
C8 phi_2 BUS[2] 0.11068f
C9 a_7084_1577# enable 0.0022f
C10 a_59860_1577# BUS[10] 0
C11 a_27432_1562# swmatrix_Tgate_5.gated_control 0.00985f
C12 a_3700_1577# enable 0.00579f
C13 a_9696_2122# a_9900_2122# 0.01151f
C14 a_9180_1580# a_9548_2122# 0.00294f
C15 a_27900_1580# phi_2 0.07395f
C16 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_23641_1539# 0.0097f
C17 a_52860_1580# BUS[9] 0.01486f
C18 a_27432_1562# phi_2 0.60119f
C19 a_59100_1580# enable 0.05124f
C20 a_52392_1562# BUS[9] 0.02518f
C21 a_58632_1562# enable 0.08694f
C22 a_18728_1562# vdd 1.00072f
C23 vdd BUS[3] 0.58892f
C24 ShiftReg_row_10_2$1_0.Q[2] a_11161_1539# 0.00241f
C25 a_7576_2002# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C26 a_3308_2122# vdd 0.00491f
C27 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C28 swmatrix_Tgate_1.gated_control a_53228_1577# 0
C29 ShiftReg_row_10_2$1_0.Q[6] a_38776_2002# 0.00242f
C30 a_19564_1577# pin 0
C31 a_16180_1577# pin 0
C32 swmatrix_Tgate_0.gated_control phi_2 0.31092f
C33 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D D_in 0.01068f
C34 a_13816_2002# swmatrix_Tgate_4.gated_control 0.01141f
C35 a_16140_2122# BUS[3] 0.00104f
C36 a_22176_2122# phi_1 0.01804f
C37 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C38 a_34508_2122# enable 0.00101f
C39 a_19712_2122# phi_1 0.01882f
C40 a_32536_2002# enable 0.05124f
C41 a_22176_2122# a_21660_1580# 0.30053f
C42 a_21192_1562# a_22176_2122# 0.07055f
C43 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45291f
C44 a_47480_2002# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C45 a_19712_2122# a_21192_1562# 0.00268f
C46 a_44156_1580# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C47 a_35000_2002# BUS[6] 0.00972f
C48 a_52860_1580# d_out 0
C49 a_31676_1580# BUS[6] 0.0049f
C50 swmatrix_Tgate_2.gated_control a_59860_1577# 0
C51 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C52 a_52392_1562# d_out 0
C53 a_37448_1562# phi_1 0.70141f
C54 ShiftReg_row_10_2$1_0.Q[8] a_50912_2122# 0.01552f
C55 a_47136_2122# a_46988_1577# 0
C56 a_45016_2002# pin 0.00117f
C57 a_844_1577# phi_2 0
C58 a_28416_2122# swmatrix_Tgate_5.gated_control 0.01553f
C59 a_7476_1577# enable 0.00577f
C60 a_28416_2122# phi_2 0.04011f
C61 a_9696_2122# a_9548_2122# 0
C62 a_9180_1580# a_10040_2002# 0.00888f
C63 a_7436_2122# enable 0.00368f
C64 a_25952_2122# swmatrix_Tgate_5.gated_control 0.01538f
C65 a_25952_2122# phi_2 0.04895f
C66 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0.00108f
C67 a_53376_2122# BUS[9] 0.01564f
C68 a_59616_2122# enable 0.11443f
C69 a_57356_2122# vdd 0.01506f
C70 a_50912_2122# BUS[9] 0.02103f
C71 pin BUS[10] 10.5929f
C72 a_57152_2122# enable 0.11055f
C73 a_6716_1580# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C74 a_3800_2002# vdd 0.32897f
C75 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C76 swmatrix_Tgate_1.gated_control a_57004_1577# 0
C77 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[4] 1.17576f
C78 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_2472_1562# 0
C79 swmatrix_Tgate_1.gated_control a_53620_1577# 0
C80 a_2472_1562# d_out 0
C81 ShiftReg_row_10_2$1_0.Q[6] a_37916_1580# 0.36203f
C82 a_37448_1562# swmatrix_Tgate_6.gated_control 0.00493f
C83 a_16280_2002# swmatrix_Tgate_4.gated_control 0.01014f
C84 a_43688_1562# phi_2 0.02762f
C85 a_12956_1580# swmatrix_Tgate_4.gated_control 0.00829f
C86 a_15788_2122# BUS[3] 0
C87 a_13816_2002# BUS[3] 0.01182f
C88 a_35000_2002# enable 0.0522f
C89 a_31676_1580# enable 0.05108f
C90 ShiftReg_row_10_2$1_0.Q[6] vdd 0.57782f
C91 a_50764_1577# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C92 swmatrix_Tgate_9.gated_control enable 0.57719f
C93 a_24968_1562# BUS[5] 0.00406f
C94 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C95 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C96 a_46620_1580# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C97 a_7084_2122# vdd 0.00491f
C98 a_46152_1562# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C99 swmatrix_Tgate_0.gated_control a_42361_1539# 0.00113f
C100 a_43688_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C101 a_34140_1580# BUS[6] 0.01486f
C102 a_54841_1539# phi_2 0
C103 a_33672_1562# BUS[6] 0.02518f
C104 a_53376_2122# d_out 0
C105 a_47480_2002# pin 0.00147f
C106 a_47136_2122# a_47380_1577# 0.01595f
C107 a_9900_2122# enable 0.00368f
C108 a_1236_1577# phi_2 0
C109 a_44156_1580# pin 0
C110 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C111 swmatrix_Tgate_2.gated_control pin 1.20655f
C112 a_9696_2122# a_10040_2002# 0.57845f
C113 a_59820_2122# vdd 0.01506f
C114 a_24968_1562# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C115 a_57004_2122# vdd 0.00491f
C116 ShiftReg_row_10_2$1_0.Q[2] a_13324_1577# 0
C117 a_28760_2002# d_out 0
C118 ShiftReg_row_10_2$1_0.Q[9] phi_1 0.05798f
C119 a_2940_1580# vdd 0.4251f
C120 a_8712_1562# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C121 swmatrix_Tgate_8.gated_control phi_1 0.01084f
C122 a_35000_2002# a_34900_1577# 0
C123 a_34140_1580# a_34508_1577# 0.00194f
C124 a_15420_1580# swmatrix_Tgate_4.gated_control 0.00668f
C125 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C126 a_16280_2002# BUS[3] 0.00972f
C127 a_14952_1562# swmatrix_Tgate_4.gated_control 0.00985f
C128 a_12956_1580# BUS[3] 0.0049f
C129 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_11161_1539# 0.0097f
C130 a_34140_1580# enable 0.05124f
C131 a_33672_1562# enable 0.08694f
C132 a_51156_1577# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C133 a_6248_1562# enable 0.08752f
C134 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C135 a_47136_2122# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C136 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_3.gated_control 0.17173f
C137 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C138 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C139 a_34656_2122# BUS[6] 0.01564f
C140 swmatrix_Tgate_0.gated_control a_40748_1577# 0
C141 a_44672_2122# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C142 a_53228_1577# phi_2 0
C143 ShiftReg_row_10_2$1_0.Q[4] a_26296_2002# 0.00242f
C144 a_32192_2122# BUS[6] 0.02103f
C145 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C146 swmatrix_Tgate_4.gated_control phi_2 0.31092f
C147 a_46620_1580# pin 0
C148 a_844_1577# D_in 0
C149 swmatrix_Tgate_3.gated_control enable 0.50853f
C150 a_3660_2122# phi_2 0.00422f
C151 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C152 a_46152_1562# pin 0.00214f
C153 a_9548_2122# enable 0.00101f
C154 a_9696_2122# a_9180_1580# 0.30053f
C155 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[9] 0.01102f
C156 a_59468_2122# vdd 0.00491f
C157 a_57496_2002# vdd 0.32602f
C158 d_out BUS[2] 0.16227f
C159 enable BUS[5] 0.21339f
C160 a_7232_2122# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C161 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C162 a_27900_1580# d_out 0
C163 a_27432_1562# d_out 0
C164 a_3456_2122# vdd 0.5594f
C165 a_34656_2122# a_34508_1577# 0
C166 ShiftReg_row_10_2$1_0.Q[6] a_38432_2122# 0.01552f
C167 a_12488_1562# phi_1 0.70141f
C168 a_20056_2002# pin 0.00117f
C169 a_15936_2122# swmatrix_Tgate_4.gated_control 0.01553f
C170 a_15420_1580# BUS[3] 0.01486f
C171 a_13472_2122# swmatrix_Tgate_4.gated_control 0.01538f
C172 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C173 a_14952_1562# BUS[3] 0.02518f
C174 a_34656_2122# enable 0.11443f
C175 a_32396_2122# vdd 0.01506f
C176 a_32192_2122# enable 0.11055f
C177 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C178 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[3] 1.17576f
C179 swmatrix_Tgate_0.gated_control d_out 0.35904f
C180 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C181 swmatrix_Tgate_0.gated_control a_44524_1577# 0
C182 swmatrix_Tgate_0.gated_control a_41140_1577# 0
C183 a_57004_1577# phi_2 0
C184 a_53620_1577# phi_2 0
C185 a_24968_1562# swmatrix_Tgate_7.gated_control 0.00493f
C186 ShiftReg_row_10_2$1_0.Q[4] a_25436_1580# 0.36203f
C187 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C188 a_18728_1562# phi_2 0.02762f
C189 a_49928_1562# enable 0.08752f
C190 phi_2 BUS[3] 0.11068f
C191 a_47136_2122# pin 0.00304f
C192 a_10040_2002# enable 0.0522f
C193 a_3308_2122# phi_2 0
C194 a_44672_2122# pin 0
C195 ShiftReg_row_10_2$1_0.Q[2] vdd 0.57782f
C196 swmatrix_Tgate_8.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00504f
C197 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0.01107f
C198 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C199 a_59960_2002# vdd 0.3289f
C200 a_56636_1580# vdd 0.42253f
C201 swmatrix_Tgate_5.gated_control a_29881_1539# 0.00113f
C202 a_31208_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C203 a_29881_1539# phi_2 0
C204 vdd BUS[4] 0.58892f
C205 a_28416_2122# d_out 0
C206 a_54841_1539# BUS[9] 0
C207 a_51116_2122# phi_1 0.00534f
C208 a_22520_2002# pin 0.00147f
C209 a_34656_2122# a_34900_1577# 0.01595f
C210 a_19196_1580# pin 0
C211 a_15936_2122# BUS[3] 0.01564f
C212 a_13472_2122# BUS[3] 0.02103f
C213 a_34860_2122# vdd 0.01506f
C214 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C215 a_32044_2122# vdd 0.00491f
C216 a_51256_2002# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C217 ShiftReg_row_10_2$1_0.Q[5] phi_1 0.05798f
C218 a_22520_2002# a_22420_1577# 0
C219 a_57396_1577# phi_2 0
C220 a_21660_1580# a_22028_1577# 0.00194f
C221 a_57356_2122# phi_2 0.00411f
C222 a_7576_2002# phi_1 0.01314f
C223 a_3800_2002# phi_2 0.03174f
C224 a_9180_1580# enable 0.05124f
C225 swmatrix_Tgate_9.gated_control a_992_2122# 0.01491f
C226 a_54841_1539# d_out 0
C227 a_59100_1580# vdd 0.4252f
C228 a_58632_1562# vdd 1.04286f
C229 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_6.gated_control 0.17173f
C230 swmatrix_Tgate_5.gated_control a_28268_1577# 0
C231 ShiftReg_row_10_2$1_0.Q[6] phi_2 0.63578f
C232 ShiftReg_row_10_2$1_0.Q[2] a_13816_2002# 0.00242f
C233 a_53580_2122# phi_1 0.00477f
C234 a_28268_1577# phi_2 0
C235 phi_1 pin 0.009f
C236 a_50764_2122# phi_1 0.00201f
C237 a_53228_1577# BUS[9] 0
C238 swmatrix_Tgate_1.gated_control a_56636_1580# 0
C239 a_56168_1562# a_57496_2002# 0.02403f
C240 swmatrix_Tgate_7.gated_control enable 0.50853f
C241 a_21660_1580# pin 0
C242 a_7084_2122# phi_2 0
C243 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C244 a_21192_1562# pin 0.00214f
C245 a_8_1562# phi_1 0.70228f
C246 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[7] 0.01102f
C247 a_53720_2002# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C248 a_34508_2122# vdd 0.00491f
C249 a_32536_2002# vdd 0.32602f
C250 a_50396_1580# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C251 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C252 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C253 a_59820_2122# phi_2 0.00422f
C254 swmatrix_Tgate_6.gated_control pin 1.20655f
C255 a_22176_2122# a_22028_1577# 0
C256 a_57004_2122# phi_2 0
C257 ShiftReg_row_10_2$1_0.Q[4] a_25952_2122# 0.01552f
C258 a_3800_2002# ShiftReg_row_10_2$1_0.Q[1] 0.25874f
C259 a_6716_1580# phi_1 0.0533f
C260 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[2] 1.17576f
C261 a_36121_1539# BUS[6] 0
C262 a_2940_1580# phi_2 0.07395f
C263 a_9696_2122# enable 0.11443f
C264 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C265 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0.08805f
C266 a_7436_2122# vdd 0.01506f
C267 a_53228_1577# d_out 0
C268 swmatrix_Tgate_4.gated_control d_out 0.35904f
C269 a_59616_2122# vdd 0.56003f
C270 a_57152_2122# vdd 0.56061f
C271 swmatrix_Tgate_3.gated_control BUS[7] 0.00677f
C272 swmatrix_Tgate_5.gated_control a_32044_1577# 0
C273 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C274 ShiftReg_row_10_2$1_0.Q[2] a_12956_1580# 0.36203f
C275 a_12488_1562# swmatrix_Tgate_8.gated_control 0.00493f
C276 swmatrix_Tgate_5.gated_control a_28660_1577# 0
C277 a_32044_1577# phi_2 0
C278 a_53228_2122# phi_1 0.00164f
C279 a_28660_1577# phi_2 0
C280 a_51256_2002# phi_1 0.01314f
C281 a_56168_1562# a_56636_1580# 0.30528f
C282 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C283 a_53620_1577# BUS[9] 0
C284 a_22176_2122# pin 0.00304f
C285 a_24968_1562# enable 0.08752f
C286 a_19712_2122# pin 0
C287 a_57004_1577# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C288 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C289 a_35000_2002# vdd 0.3289f
C290 swmatrix_Tgate_9.gated_control vdd 1.84425f
C291 a_52860_1580# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C292 a_31676_1580# vdd 0.42253f
C293 a_52392_1562# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C294 phi_1 BUS[1] 0.09502f
C295 swmatrix_Tgate_4.gated_control a_17401_1539# 0.00113f
C296 a_18728_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C297 ShiftReg_row_10_2$1_0.Q[1] ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C298 a_4921_1539# phi_2 0
C299 a_26156_2122# phi_1 0.00534f
C300 a_37448_1562# pin 0.00162f
C301 a_59468_2122# phi_2 0
C302 a_36121_1539# enable 0.00398f
C303 a_57496_2002# phi_2 0.03207f
C304 a_22176_2122# a_22420_1577# 0.01595f
C305 a_2940_1580# ShiftReg_row_10_2$1_0.Q[1] 0.00101f
C306 a_3456_2122# phi_2 0.04011f
C307 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45164f
C308 a_8712_1562# phi_1 0.01733f
C309 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C310 a_31208_1562# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C311 a_9900_2122# vdd 0.01506f
C312 a_34508_1577# BUS[6] 0
C313 a_53620_1577# d_out 0
C314 a_8_1562# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C315 d_out BUS[3] 0.16227f
C316 a_51256_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C317 enable BUS[6] 0.21339f
C318 a_32436_1577# phi_2 0
C319 a_9180_1580# a_9548_1577# 0.00194f
C320 a_10040_2002# a_9940_1577# 0
C321 a_53720_2002# phi_1 0.01261f
C322 swmatrix_Tgate_9.gated_control a_1336_2002# 0.01129f
C323 a_32396_2122# phi_2 0.00411f
C324 a_56168_1562# a_58632_1562# 0
C325 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[10] 0.10641f
C326 a_50396_1580# phi_1 0.0533f
C327 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C328 ShiftReg_row_10_2$1_0.Q[9] ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C329 a_57396_1577# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C330 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C331 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C332 a_29881_1539# d_out 0
C333 a_53376_2122# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C334 a_34140_1580# vdd 0.4252f
C335 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_7.gated_control 0.17173f
C336 a_33672_1562# vdd 1.04286f
C337 a_50912_2122# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C338 ShiftReg_row_10_2$1_0.Q[1] a_4921_1539# 0.00241f
C339 a_6248_1562# vdd 1.00072f
C340 ShiftReg_row_10_2$1_0.Q[2] phi_2 0.63578f
C341 swmatrix_Tgate_4.gated_control a_15788_1577# 0
C342 a_28620_2122# phi_1 0.00477f
C343 a_17401_1539# BUS[3] 0
C344 a_3308_1577# phi_2 0
C345 ShiftReg_row_10_2$1_0.Q[7] enable 0.513f
C346 a_25804_2122# phi_1 0.00201f
C347 a_476_1580# phi_1 0.05354f
C348 swmatrix_Tgate_0.gated_control a_44156_1580# 0
C349 a_34508_1577# enable 0.0022f
C350 a_59960_2002# phi_2 0.03174f
C351 a_43688_1562# a_45016_2002# 0.02403f
C352 swmatrix_Tgate_5.gated_control BUS[4] 0.00677f
C353 a_56636_1580# phi_2 0.03321f
C354 a_7576_2002# swmatrix_Tgate_8.gated_control 0.01141f
C355 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] 0.11433f
C356 phi_2 BUS[4] 0.11068f
C357 a_7232_2122# phi_1 0.01882f
C358 a_9548_2122# vdd 0.00491f
C359 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[5] 0.01102f
C360 swmatrix_Tgate_3.gated_control vdd 1.8044f
C361 a_34900_1577# BUS[6] 0
C362 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_53720_2002# 0.00242f
C363 ShiftReg_row_10_2$1_0.Q[9] pin 0.01625f
C364 a_50396_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C365 a_3800_2002# d_out 0
C366 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_2.gated_control 0.23535f
C367 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C368 swmatrix_Tgate_8.gated_control pin 1.20476f
C369 a_34860_2122# phi_2 0.00422f
C370 vdd BUS[5] 0.58892f
C371 ShiftReg_row_10_2$1_0.Q[2] a_13472_2122# 0.01552f
C372 a_9696_2122# a_9548_1577# 0
C373 a_32044_2122# phi_2 0
C374 a_52860_1580# phi_1 0.01277f
C375 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[1] 1.1759f
C376 a_56168_1562# a_57152_2122# 0.07055f
C377 a_52392_1562# phi_1 0.01733f
C378 ShiftReg_row_10_2$1_0.Q[6] d_out 0
C379 a_28268_1577# d_out 0
C380 a_34656_2122# vdd 0.56003f
C381 swmatrix_Tgate_4.gated_control a_19564_1577# 0
C382 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C383 swmatrix_Tgate_4.gated_control a_16180_1577# 0
C384 a_32192_2122# vdd 0.56061f
C385 a_7084_1577# phi_2 0
C386 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C387 a_28268_2122# phi_1 0.00164f
C388 a_3700_1577# phi_2 0
C389 a_38284_1577# enable 0.0022f
C390 a_15788_1577# BUS[3] 0
C391 a_43688_1562# a_44156_1580# 0.30528f
C392 a_34900_1577# enable 0.00579f
C393 a_2472_1562# phi_1 0.01733f
C394 a_26296_2002# phi_1 0.01314f
C395 a_59100_1580# phi_2 0.07395f
C396 a_6716_1580# swmatrix_Tgate_8.gated_control 0.00829f
C397 a_58632_1562# phi_2 0.60119f
C398 swmatrix_Tgate_4.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C399 a_49928_1562# vdd 1.00072f
C400 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C401 a_10040_2002# vdd 0.3289f
C402 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[7] 0.10641f
C403 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C404 swmatrix_Tgate_3.gated_control swmatrix_Tgate_1.gated_control 0.01259f
C405 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_52860_1580# 0.36162f
C406 a_50764_1577# pin 0
C407 a_47380_1577# pin 0
C408 a_52392_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C409 a_2940_1580# d_out 0
C410 a_34508_2122# phi_2 0
C411 a_11161_1539# enable 0.00398f
C412 a_2940_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C413 a_12488_1562# pin 0.00162f
C414 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[10] 0
C415 a_53376_2122# phi_1 0.01804f
C416 a_9696_2122# a_9940_1577# 0.01595f
C417 a_32536_2002# phi_2 0.03207f
C418 a_50912_2122# phi_1 0.01882f
C419 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C420 a_476_1580# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C421 swmatrix_Tgate_8.gated_control BUS[1] 0.00556f
C422 a_28660_1577# d_out 0
C423 a_57496_2002# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C424 ShiftReg_row_10_2$1_0.Q[1] a_7084_1577# 0
C425 a_38776_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C426 a_7476_1577# phi_2 0
C427 a_7436_2122# phi_2 0.00411f
C428 a_16180_1577# BUS[3] 0
C429 a_28760_2002# phi_1 0.01261f
C430 a_38676_1577# enable 0.00577f
C431 a_43688_1562# a_46152_1562# 0
C432 a_38636_2122# enable 0.00368f
C433 a_25436_1580# phi_1 0.0533f
C434 a_59616_2122# phi_2 0.04011f
C435 a_57152_2122# phi_2 0.04895f
C436 ShiftReg_row_10_2$1_0.Q[7] ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C437 a_8712_1562# swmatrix_Tgate_8.gated_control 0.00985f
C438 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_4921_1539# 0.0097f
C439 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C440 a_4921_1539# d_out 0
C441 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C442 a_59860_1577# pin 0
C443 a_9180_1580# vdd 0.4252f
C444 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C445 a_53720_2002# ShiftReg_row_10_2$1_0.Q[9] 0.25874f
C446 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C447 a_49928_1562# swmatrix_Tgate_1.gated_control 0.01446f
C448 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_53376_2122# 0.01536f
C449 a_1196_2122# phi_1 0.00534f
C450 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C451 ShiftReg_row_10_2$1_0.Q[3] enable 0.513f
C452 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_2.gated_control 0.33472f
C453 swmatrix_Tgate_3.gated_control BUS[8] 0.86839f
C454 a_31208_1562# a_32536_2002# 0.02403f
C455 a_9548_1577# enable 0.0022f
C456 swmatrix_Tgate_5.gated_control a_31676_1580# 0
C457 swmatrix_Tgate_9.gated_control phi_2 0.35589f
C458 a_3456_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C459 a_35000_2002# phi_2 0.03174f
C460 a_3456_2122# d_out 0
C461 a_31676_1580# phi_2 0.03321f
C462 swmatrix_Tgate_7.gated_control vdd 1.8044f
C463 a_2472_1562# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00423f
C464 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C465 a_59960_2002# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C466 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C467 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[3] 0.01102f
C468 a_56636_1580# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C469 ShiftReg_row_10_2$1_0.Q[5] pin 0.01625f
C470 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_41240_2002# 0.00242f
C471 a_37916_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C472 phi_1 BUS[2] 0.09482f
C473 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[4] 0.10641f
C474 a_9900_2122# phi_2 0.00422f
C475 a_27900_1580# phi_1 0.01277f
C476 a_27432_1562# phi_1 0.01733f
C477 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00187f
C478 a_41100_2122# enable 0.00368f
C479 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C480 a_38284_2122# enable 0.00101f
C481 a_43688_1562# a_44672_2122# 0.07055f
C482 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C483 a_7576_2002# pin 0.00117f
C484 a_7232_2122# swmatrix_Tgate_8.gated_control 0.01538f
C485 ShiftReg_row_10_2$1_0.Q[2] d_out 0
C486 a_3308_1577# d_out 0
C487 ShiftReg_row_10_2$1_0.Q[7] BUS[7] 0.0247f
C488 a_59960_2002# d_out 0.25884f
C489 a_9696_2122# vdd 0.56003f
C490 a_52860_1580# ShiftReg_row_10_2$1_0.Q[9] 0.00101f
C491 a_51256_2002# a_51156_1577# 0
C492 a_52392_1562# ShiftReg_row_10_2$1_0.Q[9] 0.00225f
C493 swmatrix_Tgate_0.gated_control phi_1 0.01084f
C494 a_50396_1580# a_50764_1577# 0.00194f
C495 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_9.gated_control 0.22418f
C496 a_57004_1577# swmatrix_Tgate_2.gated_control 0
C497 d_out BUS[4] 0.16227f
C498 enable BUS[7] 0.21339f
C499 a_51256_2002# a_51116_2122# 0.00109f
C500 a_13324_1577# enable 0.0022f
C501 a_34140_1580# phi_2 0.07395f
C502 a_9940_1577# enable 0.00579f
C503 a_31208_1562# a_31676_1580# 0.30528f
C504 a_6248_1562# phi_2 0.02762f
C505 a_33672_1562# phi_2 0.60119f
C506 a_57396_1577# BUS[10] 0
C507 a_8_1562# pin 0
C508 a_992_2122# enable 0.11086f
C509 a_57356_2122# BUS[10] 0
C510 a_24968_1562# vdd 1.00072f
C511 a_6716_1580# a_7576_2002# 0.00888f
C512 a_59100_1580# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C513 a_58632_1562# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C514 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C515 swmatrix_Tgate_6.gated_control swmatrix_Tgate_0.gated_control 0.01259f
C516 a_25804_1577# pin 0
C517 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_40380_1580# 0.36162f
C518 swmatrix_Tgate_3.gated_control phi_2 0.31092f
C519 a_39912_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C520 a_22420_1577# pin 0
C521 a_9548_2122# phi_2 0
C522 a_28416_2122# phi_1 0.01804f
C523 a_40748_2122# enable 0.00101f
C524 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C525 a_38776_2002# enable 0.05124f
C526 a_25952_2122# phi_1 0.01882f
C527 a_6716_1580# pin 0
C528 swmatrix_Tgate_5.gated_control BUS[5] 0.86839f
C529 a_37448_1562# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C530 phi_2 BUS[5] 0.11068f
C531 a_3700_1577# d_out 0
C532 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_3.gated_control 0.23535f
C533 a_59100_1580# d_out 0.00112f
C534 a_26296_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C535 a_58632_1562# d_out 0.00247f
C536 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] 0.11433f
C537 a_43688_1562# phi_1 0.70141f
C538 ShiftReg_row_10_2$1_0.Q[1] a_6248_1562# 0.16779f
C539 a_51256_2002# pin 0.00117f
C540 a_13716_1577# enable 0.00577f
C541 a_57396_1577# swmatrix_Tgate_2.gated_control 0
C542 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C543 a_34656_2122# phi_2 0.04011f
C544 vdd BUS[6] 0.58892f
C545 a_13676_2122# enable 0.00368f
C546 a_31208_1562# a_33672_1562# 0
C547 a_57356_2122# swmatrix_Tgate_2.gated_control 0
C548 ShiftReg_row_10_2$1_0.Q[5] ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C549 a_32192_2122# phi_2 0.04895f
C550 swmatrix_Tgate_9.gated_control D_in 0.17623f
C551 a_59820_2122# BUS[10] 0.00104f
C552 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C553 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C554 a_8712_1562# a_7576_2002# 0
C555 a_59616_2122# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C556 a_41240_2002# ShiftReg_row_10_2$1_0.Q[7] 0.25874f
C557 a_57152_2122# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C558 pin BUS[1] 10.5929f
C559 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C560 a_37448_1562# swmatrix_Tgate_0.gated_control 0.01446f
C561 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_40896_2122# 0.01536f
C562 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C563 a_8_1562# BUS[1] 0.00618f
C564 swmatrix_Tgate_4.gated_control a_19196_1580# 0
C565 a_18728_1562# a_20056_2002# 0.02403f
C566 a_49928_1562# phi_2 0.02762f
C567 ShiftReg_row_10_2$1_0.Q[4] BUS[4] 0.0247f
C568 a_10040_2002# phi_2 0.03174f
C569 a_844_2122# enable 0.00101f
C570 ShiftReg_row_10_2$1_0.Q[7] vdd 0.57782f
C571 a_41240_2002# enable 0.0522f
C572 a_37916_1580# enable 0.05108f
C573 a_8712_1562# pin 0.00214f
C574 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C575 a_38676_1577# BUS[7] 0
C576 vdd enable 4.23314f
C577 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_28760_2002# 0.00242f
C578 a_38636_2122# BUS[7] 0
C579 a_59616_2122# d_out 0.11457f
C580 a_25436_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C581 a_53720_2002# a_53580_2122# 0.00109f
C582 a_59820_2122# swmatrix_Tgate_2.gated_control 0
C583 a_50912_2122# a_50764_1577# 0
C584 a_53720_2002# pin 0.00147f
C585 a_50396_1580# a_50764_2122# 0.00294f
C586 a_16140_2122# enable 0.00368f
C587 a_50396_1580# pin 0
C588 a_13324_2122# enable 0.00101f
C589 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C590 a_31208_1562# a_32192_2122# 0.07055f
C591 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C592 a_59468_2122# BUS[10] 0
C593 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[7] 0
C594 a_57496_2002# BUS[10] 0.01182f
C595 a_844_1577# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C596 a_52860_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C597 a_52392_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C598 a_8712_1562# a_6716_1580# 0
C599 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.01636f
C600 a_7232_2122# a_7576_2002# 0.57845f
C601 a_35000_2002# d_out 0
C602 swmatrix_Tgate_8.gated_control BUS[2] 0.86839f
C603 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_9.gated_control 0.33472f
C604 a_40380_1580# ShiftReg_row_10_2$1_0.Q[7] 0.00101f
C605 swmatrix_Tgate_9.gated_control d_out 0.35905f
C606 a_38776_2002# a_38676_1577# 0
C607 swmatrix_Tgate_4.gated_control phi_1 0.01084f
C608 a_37916_1580# a_38284_1577# 0.00194f
C609 a_39912_1562# ShiftReg_row_10_2$1_0.Q[7] 0.00225f
C610 a_38776_2002# a_38636_2122# 0.00109f
C611 a_476_1580# pin 0
C612 a_18728_1562# a_19196_1580# 0.30528f
C613 a_3660_2122# phi_1 0.00477f
C614 a_9180_1580# phi_2 0.07395f
C615 a_1336_2002# enable 0.05124f
C616 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C617 swmatrix_Tgate_7.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C618 a_40380_1580# enable 0.05124f
C619 a_39912_1562# enable 0.08694f
C620 a_7232_2122# pin 0
C621 a_8_1562# a_476_1580# 0.30528f
C622 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C623 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_3.gated_control 0.22418f
C624 a_41100_2122# BUS[7] 0.00104f
C625 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_27900_1580# 0.36162f
C626 swmatrix_Tgate_7.gated_control swmatrix_Tgate_5.gated_control 0.01259f
C627 swmatrix_Tgate_7.gated_control phi_2 0.31092f
C628 a_27432_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C629 a_50912_2122# a_51156_1577# 0.01595f
C630 a_52860_1580# pin 0
C631 swmatrix_Tgate_1.gated_control enable 0.50853f
C632 a_50912_2122# a_51116_2122# 0.01151f
C633 a_50396_1580# a_51256_2002# 0.00888f
C634 a_15788_2122# enable 0.00101f
C635 a_52392_1562# pin 0.00214f
C636 a_13816_2002# enable 0.05124f
C637 a_57496_2002# swmatrix_Tgate_2.gated_control 0.01141f
C638 a_1236_1577# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C639 a_59960_2002# BUS[10] 0.00972f
C640 ShiftReg_row_10_2$1_0.Q[9] ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C641 a_56636_1580# BUS[10] 0.0049f
C642 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_53228_1577# 0
C643 a_53376_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C644 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_6.gated_control 0.23535f
C645 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C646 a_7232_2122# a_6716_1580# 0.30053f
C647 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_6248_1562# 0
C648 a_34140_1580# d_out 0
C649 a_13816_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C650 a_33672_1562# d_out 0
C651 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] 0.11433f
C652 a_18728_1562# phi_1 0.70141f
C653 phi_1 BUS[3] 0.09482f
C654 a_19956_1577# BUS[4] 0
C655 a_2472_1562# pin 0.00119f
C656 a_26296_2002# pin 0.00117f
C657 a_9696_2122# phi_2 0.04011f
C658 a_19916_2122# BUS[4] 0
C659 a_18728_1562# a_21192_1562# 0
C660 a_3308_2122# phi_1 0.00164f
C661 a_7084_1577# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C662 ShiftReg_row_10_2$1_0.Q[3] ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C663 a_40896_2122# enable 0.11443f
C664 a_38636_2122# vdd 0.01506f
C665 a_38432_2122# enable 0.11055f
C666 a_8_1562# a_2472_1562# 0
C667 swmatrix_Tgate_3.gated_control d_out 0.35904f
C668 ShiftReg_row_10_2$1_0.Q[8] a_49928_1562# 0.16779f
C669 a_44524_1577# swmatrix_Tgate_3.gated_control 0
C670 a_476_1580# BUS[1] 0.00718f
C671 a_40748_2122# BUS[7] 0
C672 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0
C673 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[4] 0
C674 a_28760_2002# ShiftReg_row_10_2$1_0.Q[5] 0.25874f
C675 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_28416_2122# 0.01536f
C676 a_24968_1562# swmatrix_Tgate_5.gated_control 0.01446f
C677 a_38776_2002# BUS[7] 0.01182f
C678 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C679 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C680 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C681 a_24968_1562# phi_2 0.02762f
C682 a_8_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C683 a_52860_1580# a_53228_2122# 0.00294f
C684 a_53376_2122# a_53580_2122# 0.01151f
C685 a_53376_2122# pin 0.00304f
C686 a_56168_1562# enable 0.08752f
C687 a_49928_1562# BUS[9] 0.00406f
C688 d_out BUS[5] 0.16227f
C689 a_59960_2002# swmatrix_Tgate_2.gated_control 0.01014f
C690 enable BUS[8] 0.21339f
C691 a_16280_2002# enable 0.0522f
C692 a_52392_1562# a_51256_2002# 0
C693 ShiftReg_row_10_2$1_0.Q[3] vdd 0.57782f
C694 a_50912_2122# pin 0
C695 a_50912_2122# a_50764_2122# 0
C696 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_59468_1577# 0
C697 a_12956_1580# enable 0.05108f
C698 a_56636_1580# swmatrix_Tgate_2.gated_control 0.00829f
C699 a_59100_1580# BUS[10] 0.01486f
C700 a_58632_1562# BUS[10] 0.02518f
C701 ShiftReg_row_10_2$1_0.Q[9] a_54841_1539# 0.00241f
C702 a_7232_2122# a_8712_1562# 0.00268f
C703 a_36121_1539# phi_2 0
C704 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_16280_2002# 0.00242f
C705 a_34656_2122# d_out 0
C706 a_12956_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C707 a_57356_2122# phi_1 0.00534f
C708 a_41240_2002# a_41100_2122# 0.00109f
C709 a_28760_2002# pin 0.00147f
C710 a_38432_2122# a_38284_1577# 0
C711 a_22380_2122# BUS[4] 0.00104f
C712 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C713 a_37916_1580# a_38284_2122# 0.00294f
C714 a_25436_1580# pin 0
C715 a_7476_1577# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C716 a_3800_2002# phi_1 0.01261f
C717 a_18728_1562# a_19712_2122# 0.07055f
C718 a_41100_2122# vdd 0.01506f
C719 a_38284_2122# vdd 0.00491f
C720 a_40380_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C721 a_39912_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C722 phi_2 BUS[6] 0.11068f
C723 a_10040_2002# d_out 0
C724 ShiftReg_row_10_2$1_0.Q[6] phi_1 0.05798f
C725 a_44916_1577# swmatrix_Tgate_3.gated_control 0
C726 a_2472_1562# BUS[1] 0.02658f
C727 a_44876_2122# swmatrix_Tgate_3.gated_control 0
C728 a_27900_1580# ShiftReg_row_10_2$1_0.Q[5] 0.00101f
C729 a_41240_2002# BUS[7] 0.00972f
C730 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C731 a_27432_1562# ShiftReg_row_10_2$1_0.Q[5] 0.00225f
C732 a_26296_2002# a_26196_1577# 0
C733 a_37916_1580# BUS[7] 0.0049f
C734 a_25436_1580# a_25804_1577# 0.00194f
C735 a_26296_2002# a_26156_2122# 0.00109f
C736 a_53376_2122# a_53228_2122# 0
C737 a_7576_2002# BUS[2] 0.01182f
C738 a_52860_1580# a_53720_2002# 0.00888f
C739 a_7084_2122# phi_1 0.00201f
C740 a_992_2122# a_844_2122# 0
C741 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_61081_1539# 0.0097f
C742 a_52392_1562# a_53720_2002# 0.02403f
C743 a_52392_1562# a_50396_1580# 0
C744 a_15420_1580# enable 0.05124f
C745 vdd BUS[7] 0.58892f
C746 a_50912_2122# a_51256_2002# 0.57845f
C747 a_59100_1580# swmatrix_Tgate_2.gated_control 0.00668f
C748 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_3.gated_control 0.33472f
C749 a_58632_1562# swmatrix_Tgate_2.gated_control 0.00985f
C750 a_14952_1562# enable 0.08694f
C751 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C752 a_59616_2122# BUS[10] 0.01564f
C753 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[1] 0.10814f
C754 a_57152_2122# BUS[10] 0.02103f
C755 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C756 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_6.gated_control 0.22418f
C757 a_992_2122# vdd 0.56059f
C758 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C759 ShiftReg_row_10_2$1_0.Q[7] phi_2 0.63578f
C760 swmatrix_Tgate_8.gated_control swmatrix_Tgate_4.gated_control 0.01259f
C761 a_34508_1577# phi_2 0
C762 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_15420_1580# 0.36162f
C763 a_59820_2122# phi_1 0.00477f
C764 pin BUS[2] 10.5929f
C765 a_14952_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C766 a_57004_2122# phi_1 0.00201f
C767 a_38432_2122# a_38676_1577# 0.01595f
C768 a_27900_1580# pin 0
C769 swmatrix_Tgate_5.gated_control enable 0.50853f
C770 a_38432_2122# a_38636_2122# 0.01151f
C771 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C772 a_27432_1562# pin 0.00214f
C773 a_37916_1580# a_38776_2002# 0.00888f
C774 a_2940_1580# phi_1 0.01277f
C775 phi_2 enable 1.58851f
C776 a_22028_2122# BUS[4] 0
C777 a_20056_2002# BUS[4] 0.01182f
C778 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C779 ShiftReg_row_10_2$1_0.Q[7] ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C780 a_40748_2122# vdd 0.00491f
C781 a_43688_1562# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C782 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_40748_1577# 0
C783 a_38776_2002# vdd 0.32602f
C784 a_40896_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C785 a_31208_1562# BUS[6] 0.00406f
C786 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_7.gated_control 0.23535f
C787 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C788 a_47340_2122# swmatrix_Tgate_3.gated_control 0
C789 a_9180_1580# d_out 0
C790 swmatrix_Tgate_0.gated_control pin 1.20655f
C791 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C792 a_40380_1580# BUS[7] 0.01486f
C793 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] 0.11433f
C794 a_39912_1562# BUS[7] 0.02518f
C795 a_6716_1580# BUS[2] 0.0049f
C796 a_992_2122# a_1336_2002# 0.57845f
C797 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C798 a_53376_2122# a_53720_2002# 0.57845f
C799 a_2472_1562# a_476_1580# 0
C800 a_59616_2122# swmatrix_Tgate_2.gated_control 0.01553f
C801 a_52392_1562# a_52860_1580# 0.30528f
C802 a_15936_2122# enable 0.11443f
C803 a_50912_2122# a_50396_1580# 0.30053f
C804 a_57152_2122# swmatrix_Tgate_2.gated_control 0.01538f
C805 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C806 a_13472_2122# enable 0.11055f
C807 a_1196_2122# BUS[1] 0.00101f
C808 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_49928_1562# 0
C809 ShiftReg_row_10_2$1_0.Q[9] a_57004_1577# 0
C810 a_13676_2122# vdd 0.01506f
C811 swmatrix_Tgate_7.gated_control d_out 0.35904f
C812 a_6248_1562# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C813 a_32044_1577# swmatrix_Tgate_6.gated_control 0
C814 a_3800_2002# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00149f
C815 ShiftReg_row_10_2$1_0.Q[6] a_37448_1562# 0.16779f
C816 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C817 a_16280_2002# ShiftReg_row_10_2$1_0.Q[3] 0.25874f
C818 a_476_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C819 a_12488_1562# swmatrix_Tgate_4.gated_control 0.01446f
C820 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_15936_2122# 0.01536f
C821 a_38284_1577# phi_2 0
C822 a_59468_2122# phi_1 0.00164f
C823 a_34900_1577# phi_2 0
C824 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C825 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C826 a_40380_1580# a_40748_2122# 0.00294f
C827 a_57496_2002# phi_1 0.01314f
C828 a_40896_2122# a_41100_2122# 0.01151f
C829 a_28416_2122# pin 0.00304f
C830 a_31208_1562# enable 0.08752f
C831 ShiftReg_row_10_2$1_0.Q[1] enable 0.513f
C832 a_38432_2122# a_38284_2122# 0
C833 a_39912_1562# a_38776_2002# 0
C834 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_54841_1539# 0.0097f
C835 a_25952_2122# pin 0
C836 a_3456_2122# phi_1 0.01804f
C837 a_22520_2002# BUS[4] 0.00972f
C838 a_19196_1580# BUS[4] 0.0049f
C839 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C840 a_844_2122# vdd 0.00491f
C841 ShiftReg_row_10_2$1_0.Q[7] a_42361_1539# 0.00241f
C842 a_41240_2002# vdd 0.3289f
C843 a_37916_1580# vdd 0.42253f
C844 a_11161_1539# phi_2 0
C845 a_32396_2122# phi_1 0.00534f
C846 a_9696_2122# d_out 0
C847 a_40896_2122# BUS[7] 0.01564f
C848 a_28760_2002# a_28620_2122# 0.00109f
C849 a_45016_2002# swmatrix_Tgate_3.gated_control 0.01141f
C850 a_42361_1539# enable 0.00398f
C851 a_43688_1562# pin 0.00162f
C852 a_25952_2122# a_25804_1577# 0
C853 a_38432_2122# BUS[7] 0.02103f
C854 a_53376_2122# a_52860_1580# 0.30053f
C855 a_25436_1580# a_25804_2122# 0.00294f
C856 a_52392_1562# a_53376_2122# 0.07055f
C857 a_8712_1562# BUS[2] 0.02518f
C858 a_50912_2122# a_52392_1562# 0.00268f
C859 a_16140_2122# vdd 0.01506f
C860 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C861 a_13324_2122# vdd 0.00491f
C862 a_27900_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C863 a_2940_1580# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00132f
C864 a_27432_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C865 a_32436_1577# swmatrix_Tgate_6.gated_control 0
C866 ShiftReg_row_10_2$1_0.Q[2] phi_1 0.05798f
C867 a_38676_1577# phi_2 0
C868 a_2472_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C869 a_32396_2122# swmatrix_Tgate_6.gated_control 0
C870 a_15420_1580# ShiftReg_row_10_2$1_0.Q[3] 0.00101f
C871 a_14952_1562# ShiftReg_row_10_2$1_0.Q[3] 0.00225f
C872 a_38636_2122# phi_2 0.00411f
C873 a_13816_2002# a_13716_1577# 0
C874 a_12956_1580# a_13324_1577# 0.00194f
C875 a_12488_1562# BUS[3] 0.00406f
C876 a_59960_2002# phi_1 0.01261f
C877 a_1236_1577# pin 0
C878 a_13816_2002# a_13676_2122# 0.00109f
C879 a_56636_1580# phi_1 0.0533f
C880 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C881 a_40896_2122# a_40748_2122# 0
C882 a_40380_1580# a_41240_2002# 0.00888f
C883 a_39912_1562# a_41240_2002# 0.02403f
C884 phi_1 BUS[4] 0.09482f
C885 a_39912_1562# a_37916_1580# 0
C886 a_21660_1580# BUS[4] 0.01486f
C887 swmatrix_Tgate_5.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C888 a_38432_2122# a_38776_2002# 0.57845f
C889 D_in enable 0.13405f
C890 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_6.gated_control 0.33472f
C891 a_21192_1562# BUS[4] 0.02518f
C892 a_10040_2002# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C893 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C894 a_36121_1539# d_out 0
C895 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C896 a_1336_2002# vdd 0.32602f
C897 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_7.gated_control 0.22418f
C898 a_40380_1580# vdd 0.4252f
C899 a_39912_1562# vdd 1.04286f
C900 a_844_1577# BUS[1] 0
C901 ShiftReg_row_10_2$1_0.Q[3] phi_2 0.63578f
C902 a_9548_1577# phi_2 0
C903 a_47480_2002# swmatrix_Tgate_3.gated_control 0.01014f
C904 ShiftReg_row_10_2$1_0.Q[8] enable 0.513f
C905 a_34860_2122# phi_1 0.00477f
C906 a_40748_1577# enable 0.0022f
C907 a_44156_1580# swmatrix_Tgate_3.gated_control 0.00829f
C908 a_32044_2122# phi_1 0.00201f
C909 a_25952_2122# a_26196_1577# 0.01595f
C910 a_25952_2122# a_26156_2122# 0.01151f
C911 a_25436_1580# a_26296_2002# 0.00888f
C912 a_7232_2122# BUS[2] 0.02103f
C913 d_out BUS[6] 0.16227f
C914 swmatrix_Tgate_1.gated_control vdd 1.8044f
C915 enable BUS[9] 0.21339f
C916 ShiftReg_row_10_2$1_0.Q[5] ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C917 a_15788_2122# vdd 0.00491f
C918 a_13816_2002# vdd 0.32602f
C919 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_28268_1577# 0
C920 a_28416_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C921 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_8.gated_control 0.23535f
C922 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C923 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C924 a_3456_2122# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00474f
C925 a_34860_2122# swmatrix_Tgate_6.gated_control 0
C926 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C927 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] 0.11433f
C928 swmatrix_Tgate_4.gated_control pin 1.20655f
C929 a_41100_2122# phi_2 0.00422f
C930 a_59100_1580# phi_1 0.01277f
C931 a_38284_2122# phi_2 0
C932 a_58632_1562# phi_1 0.01733f
C933 a_40896_2122# a_41240_2002# 0.57845f
C934 a_13324_1577# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C935 a_39912_1562# a_40380_1580# 0.30528f
C936 a_38432_2122# a_37916_1580# 0.30053f
C937 a_22176_2122# BUS[4] 0.01564f
C938 ShiftReg_row_10_2$1_0.Q[7] d_out 0
C939 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_37448_1562# 0
C940 a_9180_1580# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C941 a_19712_2122# BUS[4] 0.02103f
C942 ShiftReg_row_10_2$1_0.Q[7] a_44524_1577# 0
C943 a_34508_1577# d_out 0
C944 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C945 ShiftReg_row_10_2$1_0.Q[4] a_24968_1562# 0.16779f
C946 a_40896_2122# vdd 0.56003f
C947 a_19564_1577# swmatrix_Tgate_7.gated_control 0
C948 a_1236_1577# BUS[1] 0
C949 a_38432_2122# vdd 0.56061f
C950 phi_2 BUS[7] 0.11068f
C951 a_13324_1577# phi_2 0
C952 enable d_out 1.24595f
C953 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C954 a_44524_1577# enable 0.0022f
C955 a_34508_2122# phi_1 0.00164f
C956 a_9940_1577# phi_2 0
C957 a_46620_1580# swmatrix_Tgate_3.gated_control 0.00668f
C958 a_28416_2122# a_28620_2122# 0.01151f
C959 a_27900_1580# a_28268_2122# 0.00294f
C960 a_46152_1562# swmatrix_Tgate_3.gated_control 0.00985f
C961 a_844_1577# a_476_1580# 0.00194f
C962 a_41140_1577# enable 0.00579f
C963 a_32536_2002# phi_1 0.01314f
C964 a_25952_2122# a_25804_2122# 0
C965 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_42361_1539# 0.0097f
C966 a_27432_1562# a_26296_2002# 0
C967 a_992_2122# phi_2 0.04895f
C968 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C969 a_56168_1562# vdd 1.00072f
C970 vdd BUS[8] 0.58892f
C971 a_16280_2002# vdd 0.3289f
C972 ShiftReg_row_10_2$1_0.Q[5] a_29881_1539# 0.00241f
C973 a_12956_1580# vdd 0.42253f
C974 ShiftReg_row_10_2$1_0.Q[9] a_57496_2002# 0.00242f
C975 a_57004_1577# pin 0
C976 a_7436_2122# phi_1 0.00534f
C977 a_53620_1577# pin 0
C978 a_32536_2002# swmatrix_Tgate_6.gated_control 0.01141f
C979 a_16280_2002# a_16140_2122# 0.00109f
C980 a_40748_2122# phi_2 0
C981 a_13472_2122# a_13324_1577# 0
C982 a_17401_1539# enable 0.00398f
C983 a_18728_1562# pin 0.00162f
C984 pin BUS[3] 10.5929f
C985 a_12956_1580# a_13324_2122# 0.00294f
C986 a_59616_2122# phi_1 0.01804f
C987 a_38776_2002# phi_2 0.03207f
C988 a_57152_2122# phi_1 0.01882f
C989 a_40896_2122# a_40380_1580# 0.30053f
C990 a_13716_1577# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C991 a_39912_1562# a_40896_2122# 0.07055f
C992 a_38432_2122# a_39912_1562# 0.00268f
C993 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C994 a_15420_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C995 a_9696_2122# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C996 a_34900_1577# d_out 0
C997 a_14952_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C998 a_19956_1577# swmatrix_Tgate_7.gated_control 0
C999 a_3660_2122# BUS[1] 0.00101f
C1000 a_13716_1577# phi_2 0
C1001 a_19916_2122# swmatrix_Tgate_7.gated_control 0
C1002 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1003 a_13676_2122# phi_2 0.00411f
C1004 swmatrix_Tgate_9.gated_control phi_1 0.01701f
C1005 a_44916_1577# enable 0.00577f
C1006 a_47136_2122# swmatrix_Tgate_3.gated_control 0.01553f
C1007 a_35000_2002# phi_1 0.01261f
C1008 a_28416_2122# a_28268_2122# 0
C1009 a_27900_1580# a_28760_2002# 0.00888f
C1010 a_44876_2122# enable 0.00368f
C1011 a_31676_1580# phi_1 0.0533f
C1012 a_44672_2122# swmatrix_Tgate_3.gated_control 0.01538f
C1013 a_27432_1562# a_28760_2002# 0.02403f
C1014 a_25952_2122# a_26296_2002# 0.57845f
C1015 a_27432_1562# a_25436_1580# 0
C1016 a_11161_1539# d_out 0
C1017 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_7.gated_control 0.33472f
C1018 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C1019 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_8.gated_control 0.22418f
C1020 a_42361_1539# BUS[7] 0
C1021 a_15420_1580# vdd 0.4252f
C1022 a_14952_1562# vdd 1.04286f
C1023 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C1024 ShiftReg_row_10_2$1_0.Q[9] a_56636_1580# 0.36203f
C1025 a_56168_1562# swmatrix_Tgate_1.gated_control 0.00493f
C1026 a_844_2122# phi_2 0
C1027 a_35000_2002# swmatrix_Tgate_6.gated_control 0.01014f
C1028 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C1029 swmatrix_Tgate_1.gated_control BUS[8] 0.00677f
C1030 ShiftReg_row_10_2$1_0.Q[4] enable 0.513f
C1031 a_9900_2122# phi_1 0.00477f
C1032 a_15788_1577# enable 0.0022f
C1033 a_31676_1580# swmatrix_Tgate_6.gated_control 0.00829f
C1034 a_41240_2002# phi_2 0.03174f
C1035 a_13472_2122# a_13716_1577# 0.01595f
C1036 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C1037 a_12956_1580# a_13816_2002# 0.00888f
C1038 a_13472_2122# a_13676_2122# 0.01151f
C1039 a_37916_1580# phi_2 0.03321f
C1040 a_3800_2002# pin 0
C1041 swmatrix_Tgate_5.gated_control vdd 1.8044f
C1042 a_49928_1562# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1043 ShiftReg_row_10_2$1_0.Q[3] ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C1044 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_15788_1577# 0
C1045 vdd phi_2 4.9056f
C1046 a_15936_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C1047 ShiftReg_row_10_2$1_0.Q[6] pin 0.01625f
C1048 a_22380_2122# swmatrix_Tgate_7.gated_control 0
C1049 a_3308_2122# BUS[1] 0
C1050 a_16140_2122# phi_2 0.00422f
C1051 a_7576_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C1052 a_34140_1580# phi_1 0.01277f
C1053 a_13324_2122# phi_2 0
C1054 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1055 a_6248_1562# phi_1 0.70141f
C1056 a_33672_1562# phi_1 0.01733f
C1057 a_47340_2122# enable 0.00368f
C1058 a_28416_2122# a_28760_2002# 0.57845f
C1059 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C1060 a_27432_1562# a_27900_1580# 0.30528f
C1061 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C1062 a_44524_2122# enable 0.00101f
C1063 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C1064 a_992_2122# D_in 0.01538f
C1065 a_25952_2122# a_25436_1580# 0.30053f
C1066 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C1067 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_24968_1562# 0
C1068 ShiftReg_row_10_2$1_0.Q[3] d_out 0
C1069 ShiftReg_row_10_2$1_0.Q[5] a_32044_1577# 0
C1070 a_9548_1577# d_out 0
C1071 a_15936_2122# vdd 0.56003f
C1072 a_40748_1577# BUS[7] 0
C1073 a_13472_2122# vdd 0.56061f
C1074 ShiftReg_row_10_2$1_0.Q[2] a_12488_1562# 0.16779f
C1075 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C1076 a_7084_1577# swmatrix_Tgate_8.gated_control 0
C1077 swmatrix_Tgate_3.gated_control phi_1 0.01084f
C1078 a_52860_1580# a_53228_1577# 0.00194f
C1079 a_53720_2002# a_53620_1577# 0
C1080 a_9548_2122# phi_1 0.00164f
C1081 a_19564_1577# enable 0.0022f
C1082 a_1336_2002# phi_2 0.03207f
C1083 a_34140_1580# swmatrix_Tgate_6.gated_control 0.00668f
C1084 a_33672_1562# swmatrix_Tgate_6.gated_control 0.00985f
C1085 a_16180_1577# enable 0.00579f
C1086 a_40380_1580# phi_2 0.07395f
C1087 a_15420_1580# a_15788_2122# 0.00294f
C1088 a_15936_2122# a_16140_2122# 0.01151f
C1089 a_39912_1562# phi_2 0.60119f
C1090 a_14952_1562# a_13816_2002# 0
C1091 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_29881_1539# 0.0097f
C1092 a_2940_1580# pin 0.00124f
C1093 a_13472_2122# a_13324_2122# 0
C1094 a_6716_1580# a_7084_2122# 0.00294f
C1095 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C1096 phi_1 BUS[5] 0.09482f
C1097 a_31208_1562# vdd 1.00072f
C1098 a_13816_2002# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1099 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C1100 ShiftReg_row_10_2$1_0.Q[1] vdd 0.57798f
C1101 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C1102 ShiftReg_row_10_2$1_0.Q[3] a_17401_1539# 0.00241f
C1103 ShiftReg_row_10_2$1_0.Q[7] a_45016_2002# 0.00242f
C1104 a_32044_1577# pin 0
C1105 a_28660_1577# pin 0
C1106 a_3800_2002# BUS[1] 0.01083f
C1107 a_20056_2002# swmatrix_Tgate_7.gated_control 0.01141f
C1108 swmatrix_Tgate_1.gated_control phi_2 0.31092f
C1109 a_6716_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C1110 a_15788_2122# phi_2 0
C1111 a_23641_1539# BUS[4] 0
C1112 a_46988_2122# enable 0.00101f
C1113 a_34656_2122# phi_1 0.01804f
C1114 a_13816_2002# phi_2 0.03207f
C1115 a_28416_2122# a_27900_1580# 0.30053f
C1116 a_32192_2122# phi_1 0.01882f
C1117 a_45016_2002# enable 0.05124f
C1118 a_27432_1562# a_28416_2122# 0.07055f
C1119 swmatrix_Tgate_6.gated_control BUS[5] 0.00677f
C1120 a_25952_2122# a_27432_1562# 0.00268f
C1121 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C1122 d_out BUS[7] 0.16227f
C1123 a_9940_1577# d_out 0
C1124 enable BUS[10] 0.21339f
C1125 a_59100_1580# a_59468_1577# 0.00194f
C1126 a_59960_2002# a_59860_1577# 0
C1127 a_41140_1577# BUS[7] 0
C1128 a_7476_1577# swmatrix_Tgate_8.gated_control 0
C1129 a_49928_1562# phi_1 0.70141f
C1130 a_7436_2122# swmatrix_Tgate_8.gated_control 0
C1131 ShiftReg_row_10_2$1_0.Q[9] a_57152_2122# 0.01552f
C1132 a_10040_2002# phi_1 0.01261f
C1133 a_53376_2122# a_53228_1577# 0
C1134 a_34656_2122# swmatrix_Tgate_6.gated_control 0.01553f
C1135 a_57496_2002# pin 0.00117f
C1136 a_19956_1577# enable 0.00577f
C1137 a_19916_2122# enable 0.00368f
C1138 a_15936_2122# a_15788_2122# 0
C1139 a_40896_2122# phi_2 0.04011f
C1140 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C1141 a_32192_2122# swmatrix_Tgate_6.gated_control 0.01538f
C1142 a_15420_1580# a_16280_2002# 0.00888f
C1143 a_14952_1562# a_16280_2002# 0.02403f
C1144 a_38432_2122# phi_2 0.04895f
C1145 a_3456_2122# pin 0.00232f
C1146 swmatrix_Tgate_6.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C1147 a_13472_2122# a_13816_2002# 0.57845f
C1148 a_14952_1562# a_12956_1580# 0
C1149 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_8.gated_control 0.33472f
C1150 a_16280_2002# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C1151 a_12956_1580# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1152 vdd D_in 0.18929f
C1153 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C1154 a_43688_1562# swmatrix_Tgate_0.gated_control 0.00493f
C1155 ShiftReg_row_10_2$1_0.Q[7] a_44156_1580# 0.36203f
C1156 a_56168_1562# phi_2 0.02762f
C1157 a_22520_2002# swmatrix_Tgate_7.gated_control 0.01014f
C1158 a_19196_1580# swmatrix_Tgate_7.gated_control 0.00829f
C1159 phi_2 BUS[8] 0.11068f
C1160 a_2940_1580# BUS[1] 0.01275f
C1161 a_16280_2002# phi_2 0.03174f
C1162 swmatrix_Tgate_9.gated_control swmatrix_Tgate_8.gated_control 0.01259f
C1163 a_8712_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C1164 a_12956_1580# phi_2 0.03321f
C1165 a_22028_1577# BUS[4] 0
C1166 ShiftReg_row_10_2$1_0.Q[8] vdd 0.57782f
C1167 a_47480_2002# enable 0.0522f
C1168 a_44156_1580# enable 0.05108f
C1169 swmatrix_Tgate_2.gated_control enable 0.50439f
C1170 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C1171 a_59616_2122# a_59468_1577# 0
C1172 a_49928_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C1173 vdd BUS[9] 0.58892f
C1174 swmatrix_Tgate_3.gated_control a_48601_1539# 0.00113f
C1175 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[8] 0.10641f
C1176 ShiftReg_row_10_2$1_0.Q[2] pin 0.01625f
C1177 a_9900_2122# swmatrix_Tgate_8.gated_control 0
C1178 a_53376_2122# a_53620_1577# 0.01595f
C1179 a_59960_2002# pin 0.00147f
C1180 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98523f
C1181 a_56636_1580# pin 0
C1182 a_1336_2002# D_in 0.00242f
C1183 a_22380_2122# enable 0.00368f
C1184 a_9180_1580# phi_1 0.01277f
C1185 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C1186 a_15936_2122# a_16280_2002# 0.57845f
C1187 a_19564_2122# enable 0.00101f
C1188 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C1189 a_14952_1562# a_15420_1580# 0.30528f
C1190 pin BUS[4] 10.5929f
C1191 a_19564_1577# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1192 a_13472_2122# a_12956_1580# 0.30053f
C1193 a_4921_1539# BUS[1] 0
C1194 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_12488_1562# 0
C1195 a_7232_2122# a_7084_2122# 0
C1196 ShiftReg_row_10_2$1_0.Q[3] a_19564_1577# 0
C1197 a_15420_1580# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C1198 a_14952_1562# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C1199 a_41240_2002# d_out 0
C1200 swmatrix_Tgate_4.gated_control BUS[2] 0.00677f
C1201 a_40380_1580# a_40748_1577# 0.00194f
C1202 swmatrix_Tgate_7.gated_control phi_1 0.01084f
C1203 a_41240_2002# a_41140_1577# 0
C1204 a_6248_1562# swmatrix_Tgate_8.gated_control 0.01446f
C1205 a_21660_1580# swmatrix_Tgate_7.gated_control 0.00668f
C1206 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1207 a_15420_1580# phi_2 0.07395f
C1208 a_3456_2122# BUS[1] 0.01544f
C1209 a_22420_1577# BUS[4] 0
C1210 a_21192_1562# swmatrix_Tgate_7.gated_control 0.00985f
C1211 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.42832f
C1212 a_14952_1562# phi_2 0.60119f
C1213 vdd d_out 20.7282f
C1214 a_46620_1580# enable 0.05124f
C1215 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_17401_1539# 0.0097f
C1216 a_3800_2002# a_2472_1562# 0.02403f
C1217 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C1218 a_46152_1562# enable 0.08694f
C1219 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_1.gated_control 0.17173f
C1220 swmatrix_Tgate_3.gated_control a_46988_1577# 0
C1221 a_59616_2122# a_59860_1577# 0.01595f
C1222 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C1223 a_7084_1577# pin 0
C1224 ShiftReg_row_10_2$1_0.Q[5] a_32536_2002# 0.00242f
C1225 a_3700_1577# pin 0
C1226 swmatrix_Tgate_5.gated_control phi_2 0.31092f
C1227 a_3800_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00242f
C1228 swmatrix_Tgate_1.gated_control BUS[9] 0.86839f
C1229 a_59100_1580# pin 0
C1230 a_9696_2122# phi_1 0.01804f
C1231 a_58632_1562# pin 0.00214f
C1232 a_22028_2122# enable 0.00101f
C1233 a_20056_2002# enable 0.05124f
C1234 a_19956_1577# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1235 a_15936_2122# a_15420_1580# 0.30053f
C1236 a_14952_1562# a_15936_2122# 0.07055f
C1237 a_13472_2122# a_14952_1562# 0.00268f
C1238 a_15936_2122# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C1239 a_3308_1577# BUS[1] 0
C1240 a_13472_2122# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1241 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C1242 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C1243 a_40380_1580# d_out 0
C1244 a_39912_1562# d_out 0
C1245 a_24968_1562# phi_1 0.70141f
C1246 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1247 ShiftReg_row_10_2$1_0.Q[7] a_44672_2122# 0.01552f
C1248 a_40896_2122# a_40748_1577# 0
C1249 a_7576_2002# a_7476_1577# 0
C1250 a_8712_1562# ShiftReg_row_10_2$1_0.Q[2] 0.00225f
C1251 a_22176_2122# swmatrix_Tgate_7.gated_control 0.01553f
C1252 a_6716_1580# a_7084_1577# 0.00194f
C1253 a_32536_2002# pin 0.00117f
C1254 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[5] 0.10641f
C1255 a_19712_2122# swmatrix_Tgate_7.gated_control 0.01538f
C1256 a_15936_2122# phi_2 0.04011f
C1257 a_7576_2002# a_7436_2122# 0.00109f
C1258 a_13472_2122# phi_2 0.04895f
C1259 a_47136_2122# enable 0.11443f
C1260 a_2940_1580# a_2472_1562# 0.30528f
C1261 a_44672_2122# enable 0.11055f
C1262 a_44876_2122# vdd 0.01506f
C1263 swmatrix_Tgate_1.gated_control d_out 0.35904f
C1264 swmatrix_Tgate_3.gated_control a_50764_1577# 0
C1265 ShiftReg_row_10_2$1_0.Q[8] BUS[8] 0.0247f
C1266 swmatrix_Tgate_3.gated_control a_47380_1577# 0
C1267 ShiftReg_row_10_2$1_0.Q[5] a_31676_1580# 0.36203f
C1268 a_31208_1562# swmatrix_Tgate_5.gated_control 0.00493f
C1269 a_10040_2002# swmatrix_Tgate_8.gated_control 0.01014f
C1270 ShiftReg_row_10_2$1_0.Q[1] phi_2 0.63578f
C1271 a_31208_1562# phi_2 0.02762f
C1272 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C1273 a_2940_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.36162f
C1274 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C1275 a_59616_2122# pin 0.00304f
C1276 a_57152_2122# pin 0
C1277 a_22520_2002# enable 0.0522f
C1278 ShiftReg_row_10_2$1_0.Q[4] vdd 0.57782f
C1279 a_19196_1580# enable 0.05108f
C1280 a_56168_1562# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1281 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C1282 a_3700_1577# BUS[1] 0
C1283 phi_1 BUS[6] 0.09482f
C1284 swmatrix_Tgate_6.gated_control a_36121_1539# 0.00113f
C1285 a_37448_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C1286 a_42361_1539# phi_2 0
C1287 a_40896_2122# d_out 0
C1288 a_35000_2002# pin 0.00147f
C1289 a_40896_2122# a_41140_1577# 0.01595f
C1290 swmatrix_Tgate_9.gated_control pin 1.18579f
C1291 a_31676_1580# pin 0
C1292 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1293 a_47340_2122# vdd 0.01506f
C1294 swmatrix_Tgate_9.gated_control a_8_1562# 0.01228f
C1295 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C1296 a_44524_2122# vdd 0.00491f
C1297 a_3456_2122# a_2472_1562# 0.07055f
C1298 swmatrix_Tgate_6.gated_control BUS[6] 0.86839f
C1299 d_out BUS[8] 0.16227f
C1300 ShiftReg_row_10_2$1_0.Q[7] phi_1 0.05798f
C1301 a_16280_2002# d_out 0
C1302 a_27900_1580# a_28268_1577# 0.00194f
C1303 a_28760_2002# a_28660_1577# 0
C1304 a_9180_1580# swmatrix_Tgate_8.gated_control 0.00668f
C1305 D_in phi_2 0.36302f
C1306 a_3456_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01536f
C1307 phi_1 enable 0.69314f
C1308 a_21660_1580# enable 0.05124f
C1309 swmatrix_Tgate_9.gated_control a_6716_1580# 0
C1310 a_6248_1562# a_7576_2002# 0.02403f
C1311 a_21192_1562# enable 0.08694f
C1312 a_20056_2002# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1313 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[2] 0.10641f
C1314 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_0.gated_control 0.17173f
C1315 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C1316 swmatrix_Tgate_6.gated_control a_34508_1577# 0
C1317 ShiftReg_row_10_2$1_0.Q[3] a_20056_2002# 0.00242f
C1318 ShiftReg_row_10_2$1_0.Q[8] phi_2 0.63578f
C1319 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98611f
C1320 a_40748_1577# phi_2 0
C1321 swmatrix_Tgate_6.gated_control enable 0.50853f
C1322 a_34140_1580# pin 0
C1323 ShiftReg_row_10_2$1_0.Q[5] BUS[5] 0.0247f
C1324 a_6248_1562# pin 0.00162f
C1325 phi_2 BUS[9] 0.11068f
C1326 a_33672_1562# pin 0.00214f
C1327 a_7232_2122# a_7084_1577# 0
C1328 a_46988_2122# vdd 0.00491f
C1329 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[8] 0.01102f
C1330 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C1331 a_45016_2002# vdd 0.32602f
C1332 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_3308_1577# 0
C1333 swmatrix_Tgate_9.gated_control BUS[1] 0.86839f
C1334 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C1335 a_8712_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1336 a_44916_1577# BUS[8] 0
C1337 vdd BUS[10] 0.58892f
C1338 a_15420_1580# d_out 0
C1339 a_14952_1562# d_out 0
C1340 swmatrix_Tgate_3.gated_control pin 1.20655f
C1341 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C1342 a_44876_2122# BUS[8] 0
C1343 a_28416_2122# a_28268_1577# 0
C1344 ShiftReg_row_10_2$1_0.Q[5] a_32192_2122# 0.01552f
C1345 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C1346 a_9696_2122# swmatrix_Tgate_8.gated_control 0.01553f
C1347 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C1348 swmatrix_Tgate_0.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C1349 a_22176_2122# enable 0.11443f
C1350 pin BUS[5] 10.5929f
C1351 a_6248_1562# a_6716_1580# 0.30528f
C1352 a_19712_2122# enable 0.11055f
C1353 a_19916_2122# vdd 0.01506f
C1354 a_22520_2002# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C1355 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[8] 0
C1356 swmatrix_Tgate_5.gated_control d_out 0.35904f
C1357 a_19196_1580# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1358 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C1359 swmatrix_Tgate_6.gated_control a_38284_1577# 0
C1360 phi_2 d_out 0.66837f
C1361 a_44524_1577# phi_2 0
C1362 swmatrix_Tgate_6.gated_control a_34900_1577# 0
C1363 a_18728_1562# swmatrix_Tgate_4.gated_control 0.00493f
C1364 ShiftReg_row_10_2$1_0.Q[3] a_19196_1580# 0.36203f
C1365 a_41140_1577# phi_2 0
C1366 swmatrix_Tgate_4.gated_control BUS[3] 0.86839f
C1367 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C1368 a_34656_2122# pin 0.00304f
C1369 a_37448_1562# enable 0.08752f
C1370 a_32192_2122# pin 0
C1371 a_7232_2122# a_7476_1577# 0.01595f
C1372 a_7232_2122# a_7436_2122# 0.01151f
C1373 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C1374 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C1375 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.10961f
C1376 a_47480_2002# vdd 0.3289f
C1377 a_44156_1580# vdd 0.42253f
C1378 swmatrix_Tgate_2.gated_control vdd 1.804f
C1379 swmatrix_Tgate_7.gated_control a_23641_1539# 0.00113f
C1380 a_24968_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C1381 a_17401_1539# phi_2 0
C1382 a_15936_2122# d_out 0
C1383 a_49928_1562# pin 0.00162f
C1384 a_38636_2122# phi_1 0.00534f
C1385 a_47340_2122# BUS[8] 0.00104f
C1386 a_48601_1539# enable 0.00398f
C1387 a_28416_2122# a_28660_1577# 0.01595f
C1388 a_10040_2002# pin 0.00147f
C1389 swmatrix_Tgate_9.gated_control a_476_1580# 0.00815f
C1390 a_25804_1577# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1391 a_22380_2122# vdd 0.01506f
C1392 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C1393 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C1394 a_6248_1562# a_8712_1562# 0
C1395 a_19564_2122# vdd 0.00491f
C1396 a_21660_1580# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C1397 ShiftReg_row_10_2$1_0.Q[1] ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C1398 a_21192_1562# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C1399 ShiftReg_row_10_2$1_0.Q[1] d_out 0
C1400 ShiftReg_row_10_2$1_0.Q[2] BUS[2] 0.0247f
C1401 a_57496_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C1402 ShiftReg_row_10_2$1_0.Q[3] phi_1 0.05798f
C1403 a_44916_1577# phi_2 0
C1404 a_15420_1580# a_15788_1577# 0.00194f
C1405 a_16280_2002# a_16180_1577# 0
C1406 a_44876_2122# phi_2 0.00411f
C1407 a_3800_2002# a_3660_2122# 0.00109f
C1408 a_26196_1577# BUS[5] 0
C1409 a_42361_1539# d_out 0
C1410 a_26156_2122# BUS[5] 0
C1411 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C1412 a_46620_1580# vdd 0.4252f
C1413 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_5.gated_control 0.17173f
C1414 a_61081_1539# enable 0.00398f
C1415 swmatrix_Tgate_7.gated_control a_22028_1577# 0
C1416 a_46152_1562# vdd 1.04286f
C1417 ShiftReg_row_10_2$1_0.Q[4] phi_2 0.63578f
C1418 a_41100_2122# phi_1 0.00477f
C1419 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[5] 0
C1420 ShiftReg_row_10_2$1_0.Q[9] enable 0.513f
C1421 a_15788_1577# phi_2 0
C1422 a_46988_2122# BUS[8] 0
C1423 a_46988_1577# enable 0.0022f
C1424 swmatrix_Tgate_3.gated_control a_50396_1580# 0
C1425 a_49928_1562# a_51256_2002# 0.02403f
C1426 a_38284_2122# phi_1 0.00201f
C1427 swmatrix_Tgate_8.gated_control enable 0.50853f
C1428 swmatrix_Tgate_1.gated_control swmatrix_Tgate_2.gated_control 0.01259f
C1429 a_45016_2002# BUS[8] 0.01182f
C1430 a_9180_1580# pin 0
C1431 swmatrix_Tgate_9.gated_control a_2472_1562# 0.00985f
C1432 a_56168_1562# BUS[10] 0.00406f
C1433 a_26196_1577# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1434 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[6] 0.01102f
C1435 a_22028_2122# vdd 0.00491f
C1436 a_20056_2002# vdd 0.32602f
C1437 a_22176_2122# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C1438 a_6248_1562# a_7232_2122# 0.07055f
C1439 a_19712_2122# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1440 phi_1 BUS[7] 0.09482f
C1441 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_59960_2002# 0.00242f
C1442 a_56636_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C1443 swmatrix_Tgate_9.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.23535f
C1444 a_15936_2122# a_15788_1577# 0
C1445 a_47340_2122# phi_2 0.00422f
C1446 swmatrix_Tgate_7.gated_control pin 1.20655f
C1447 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C1448 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1449 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C1450 ShiftReg_row_10_2$1_0.Q[3] a_19712_2122# 0.01552f
C1451 a_44524_2122# phi_2 0
C1452 a_992_2122# phi_1 0.01882f
C1453 a_28620_2122# BUS[5] 0.00104f
C1454 a_8712_1562# a_10040_2002# 0.02403f
C1455 ShiftReg_row_10_2$1_0.Q[8] d_out 0
C1456 a_40748_1577# d_out 0
C1457 a_47136_2122# vdd 0.56003f
C1458 a_44672_2122# vdd 0.56061f
C1459 swmatrix_Tgate_7.gated_control a_25804_1577# 0
C1460 a_59468_1577# enable 0.0022f
C1461 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C1462 swmatrix_Tgate_7.gated_control a_22420_1577# 0
C1463 a_19564_1577# phi_2 0
C1464 d_out BUS[9] 0.16227f
C1465 a_16180_1577# phi_2 0
C1466 a_50764_1577# enable 0.0022f
C1467 a_40748_2122# phi_1 0.00164f
C1468 a_47480_2002# BUS[8] 0.00972f
C1469 a_49928_1562# a_50396_1580# 0.30528f
C1470 a_44156_1580# BUS[8] 0.0049f
C1471 a_47380_1577# enable 0.00579f
C1472 a_38776_2002# phi_1 0.01314f
C1473 a_9696_2122# pin 0.00304f
C1474 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C1475 a_12488_1562# enable 0.08752f
C1476 a_56168_1562# swmatrix_Tgate_2.gated_control 0.01446f
C1477 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.47261f
C1478 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C1479 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C1480 a_22520_2002# vdd 0.3289f
C1481 swmatrix_Tgate_8.gated_control a_11161_1539# 0.00113f
C1482 a_19196_1580# vdd 0.42253f
C1483 a_12488_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C1484 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_59100_1580# 0.36162f
C1485 a_7476_1577# BUS[2] 0
C1486 a_58632_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C1487 a_7436_2122# BUS[2] 0
C1488 swmatrix_Tgate_9.gated_control a_1196_2122# 0
C1489 a_13676_2122# phi_1 0.00534f
C1490 a_24968_1562# pin 0.00162f
C1491 a_23641_1539# enable 0.00398f
C1492 a_15936_2122# a_16180_1577# 0.01595f
C1493 a_46988_2122# phi_2 0
C1494 a_45016_2002# phi_2 0.03207f
C1495 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1496 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C1497 a_28268_2122# BUS[5] 0
C1498 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[2] 0
C1499 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C1500 phi_2 BUS[10] 0.11068f
C1501 a_26296_2002# BUS[5] 0.01182f
C1502 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C1503 a_8712_1562# a_9180_1580# 0.30528f
C1504 a_3456_2122# a_3660_2122# 0.01151f
C1505 a_2940_1580# a_3308_2122# 0.00294f
C1506 a_41140_1577# d_out 0
C1507 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C1508 a_45016_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C1509 a_37448_1562# BUS[7] 0.00406f
C1510 a_59860_1577# enable 0.00579f
C1511 a_844_2122# phi_1 0.00201f
C1512 a_19956_1577# phi_2 0
C1513 a_41240_2002# phi_1 0.01261f
C1514 a_19916_2122# phi_2 0.00411f
C1515 a_51156_1577# enable 0.00577f
C1516 a_37916_1580# phi_1 0.0533f
C1517 a_46620_1580# BUS[8] 0.01486f
C1518 a_51116_2122# enable 0.00368f
C1519 a_46152_1562# BUS[8] 0.02518f
C1520 a_49928_1562# a_52392_1562# 0
C1521 ShiftReg_row_10_2$1_0.Q[8] ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C1522 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1523 a_26296_2002# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1524 a_17401_1539# d_out 0
C1525 vdd phi_1 9.99921f
C1526 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C1527 a_21660_1580# vdd 0.4252f
C1528 a_992_2122# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1529 a_21192_1562# vdd 1.04286f
C1530 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C1531 pin BUS[6] 10.5929f
C1532 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_4.gated_control 0.17173f
C1533 swmatrix_Tgate_8.gated_control a_9548_1577# 0
C1534 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_59616_2122# 0.01536f
C1535 a_9900_2122# BUS[2] 0.00104f
C1536 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1537 a_16140_2122# phi_1 0.00477f
C1538 ShiftReg_row_10_2$1_0.Q[5] enable 0.513f
C1539 a_47480_2002# phi_2 0.03174f
C1540 a_13324_2122# phi_1 0.00201f
C1541 swmatrix_Tgate_6.gated_control a_37916_1580# 0
C1542 a_22028_1577# enable 0.0022f
C1543 a_37448_1562# a_38776_2002# 0.02403f
C1544 a_44156_1580# phi_2 0.03321f
C1545 swmatrix_Tgate_2.gated_control phi_2 0.31092f
C1546 a_7576_2002# enable 0.05124f
C1547 swmatrix_Tgate_6.gated_control vdd 1.8044f
C1548 a_28760_2002# BUS[5] 0.00972f
C1549 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[4] 0.01102f
C1550 a_8712_1562# a_9696_2122# 0.07055f
C1551 a_3456_2122# a_3308_2122# 0
C1552 a_2940_1580# a_3800_2002# 0.00888f
C1553 a_25436_1580# BUS[5] 0.0049f
C1554 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_47480_2002# 0.00242f
C1555 ShiftReg_row_10_2$1_0.Q[7] pin 0.01625f
C1556 a_44156_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C1557 a_22380_2122# phi_2 0.00422f
C1558 a_1336_2002# phi_1 0.01314f
C1559 a_19564_2122# phi_2 0
C1560 a_53580_2122# enable 0.00368f
C1561 a_844_1577# swmatrix_Tgate_9.gated_control 0
C1562 a_40380_1580# phi_1 0.01277f
C1563 a_6248_1562# BUS[2] 0.00406f
C1564 a_49928_1562# a_50912_2122# 0.07055f
C1565 a_39912_1562# phi_1 0.01733f
C1566 enable pin 1.13379f
C1567 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C1568 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C1569 a_47136_2122# BUS[8] 0.01564f
C1570 a_50764_2122# enable 0.00101f
C1571 a_44672_2122# BUS[8] 0.02103f
C1572 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C1573 swmatrix_Tgate_3.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C1574 a_28760_2002# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C1575 a_8_1562# enable 0.08872f
C1576 ShiftReg_row_10_2$1_0.Q[4] d_out 0
C1577 a_25436_1580# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1578 a_15788_1577# d_out 0
C1579 a_22176_2122# vdd 0.56003f
C1580 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C1581 a_19712_2122# vdd 0.56061f
C1582 swmatrix_Tgate_8.gated_control a_13324_1577# 0
C1583 swmatrix_Tgate_8.gated_control a_9940_1577# 0
C1584 a_59100_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1585 a_9548_2122# BUS[2] 0
C1586 a_56636_1580# a_57004_1577# 0.00194f
C1587 a_58632_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1588 a_15788_2122# phi_1 0.00164f
C1589 a_57496_2002# a_57396_1577# 0
C1590 swmatrix_Tgate_1.gated_control phi_1 0.01084f
C1591 a_57496_2002# a_57356_2122# 0.00109f
C1592 a_25804_1577# enable 0.0022f
C1593 a_13816_2002# phi_1 0.01314f
C1594 a_46620_1580# phi_2 0.07395f
C1595 a_22420_1577# enable 0.00579f
C1596 a_37448_1562# a_37916_1580# 0.30528f
C1597 a_46152_1562# phi_2 0.60119f
C1598 a_18728_1562# BUS[4] 0.00406f
C1599 a_6716_1580# enable 0.05108f
C1600 a_27900_1580# BUS[5] 0.01486f
C1601 a_37448_1562# vdd 1.00072f
C1602 a_3456_2122# a_3800_2002# 0.57845f
C1603 a_27432_1562# BUS[5] 0.02518f
C1604 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_46620_1580# 0.36162f
C1605 swmatrix_Tgate_0.gated_control swmatrix_Tgate_3.gated_control 0.01259f
C1606 a_38284_1577# pin 0
C1607 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.99095f
C1608 a_46152_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C1609 a_34900_1577# pin 0
C1610 a_22028_2122# phi_2 0
C1611 a_20056_2002# phi_2 0.03207f
C1612 a_1236_1577# swmatrix_Tgate_9.gated_control 0
C1613 a_40896_2122# phi_1 0.01804f
C1614 a_53228_2122# enable 0.00101f
C1615 a_32044_1577# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1616 a_38432_2122# phi_1 0.01882f
C1617 a_51256_2002# enable 0.05124f
C1618 a_27900_1580# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C1619 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C1620 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_1.gated_control 0.23535f
C1621 a_16180_1577# d_out 0
C1622 a_27432_1562# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C1623 a_59616_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C1624 a_32536_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C1625 a_56168_1562# phi_1 0.70141f
C1626 a_10040_2002# BUS[2] 0.00972f
C1627 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[10] 1.17576f
C1628 enable BUS[1] 0.22178f
C1629 a_26196_1577# enable 0.00577f
C1630 phi_1 BUS[8] 0.09482f
C1631 a_16280_2002# phi_1 0.01261f
C1632 a_12956_1580# phi_1 0.0533f
C1633 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C1634 a_26156_2122# enable 0.00368f
C1635 a_37448_1562# a_39912_1562# 0
C1636 a_47136_2122# phi_2 0.04011f
C1637 ShiftReg_row_10_2$1_0.Q[6] ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C1638 a_44672_2122# phi_2 0.04895f
C1639 a_1336_2002# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1640 a_28416_2122# BUS[5] 0.01564f
C1641 a_8712_1562# enable 0.08694f
C1642 a_3456_2122# a_2940_1580# 0.30053f
C1643 a_25952_2122# BUS[5] 0.02103f
C1644 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C1645 a_47480_2002# ShiftReg_row_10_2$1_0.Q[8] 0.25874f
C1646 a_43688_1562# swmatrix_Tgate_3.gated_control 0.01446f
C1647 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_47136_2122# 0.01536f
C1648 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1649 a_24968_1562# a_26296_2002# 0.02403f
C1650 swmatrix_Tgate_7.gated_control a_25436_1580# 0
C1651 a_22520_2002# phi_2 0.03174f
C1652 d_out BUS[10] 0.19472f
C1653 a_19196_1580# phi_2 0.03321f
C1654 a_53720_2002# enable 0.0522f
C1655 a_3660_2122# swmatrix_Tgate_9.gated_control 0
C1656 ShiftReg_row_10_2$1_0.Q[9] vdd 0.57782f
C1657 a_50396_1580# enable 0.05108f
C1658 a_32436_1577# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1659 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C1660 swmatrix_Tgate_8.gated_control vdd 1.8009f
C1661 swmatrix_Tgate_2.gated_control BUS[9] 0.00677f
C1662 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D ShiftReg_row_10_2$1_0.Q[2] 0.01102f
C1663 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C1664 a_28416_2122# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C1665 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C1666 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_35000_2002# 0.00242f
C1667 ShiftReg_row_10_2$1_0.Q[3] pin 0.01625f
C1668 a_25952_2122# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1669 a_31676_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C1670 a_59960_2002# a_59820_2122# 0.00109f
C1671 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1672 a_57152_2122# a_57004_1577# 0
C1673 a_9180_1580# BUS[2] 0.01486f
C1674 a_15420_1580# phi_1 0.01277f
C1675 a_28620_2122# enable 0.00368f
C1676 a_56636_1580# a_57004_2122# 0.00294f
C1677 a_14952_1562# phi_1 0.01733f
C1678 a_25804_2122# enable 0.00101f
C1679 a_3800_2002# a_3700_1577# 0
C1680 a_2940_1580# a_3308_1577# 0.00194f
C1681 a_37448_1562# a_38432_2122# 0.07055f
C1682 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C1683 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C1684 a_476_1580# enable 0.05187f
C1685 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C1686 a_7232_2122# enable 0.11055f
C1687 a_47480_2002# d_out 0
C1688 a_46620_1580# ShiftReg_row_10_2$1_0.Q[8] 0.00101f
C1689 swmatrix_Tgate_2.gated_control d_out 0.59173f
C1690 swmatrix_Tgate_5.gated_control phi_1 0.01084f
C1691 a_44156_1580# a_44524_1577# 0.00194f
C1692 a_45016_2002# a_44916_1577# 0
C1693 a_46152_1562# ShiftReg_row_10_2$1_0.Q[8] 0.00225f
C1694 phi_1 phi_2 25.4284f
C1695 a_45016_2002# a_44876_2122# 0.00109f
C1696 a_24968_1562# a_25436_1580# 0.30528f
C1697 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C1698 a_21660_1580# phi_2 0.07395f
C1699 a_52860_1580# enable 0.05124f
C1700 a_21192_1562# phi_2 0.60119f
C1701 a_52392_1562# enable 0.08694f
C1702 a_12488_1562# vdd 1.00072f
C1703 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_1.gated_control 0.22418f
C1704 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C1705 pin BUS[7] 10.5929f
C1706 swmatrix_Tgate_5.gated_control swmatrix_Tgate_6.gated_control 0.01259f
C1707 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_34140_1580# 0.36162f
C1708 a_13324_1577# pin 0
C1709 a_48601_1539# BUS[8] 0
C1710 a_9940_1577# pin 0
C1711 a_33672_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C1712 swmatrix_Tgate_6.gated_control phi_2 0.31092f
C1713 a_57152_2122# a_57396_1577# 0.01595f
C1714 a_9696_2122# BUS[2] 0.01564f
C1715 a_3456_2122# a_3308_1577# 0
C1716 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1717 a_15936_2122# phi_1 0.01804f
C1718 a_56636_1580# a_57496_2002# 0.00888f
C1719 a_28268_2122# enable 0.00101f
C1720 a_992_2122# pin 0.00146f
C1721 a_57152_2122# a_57356_2122# 0.01151f
C1722 a_13472_2122# phi_1 0.01882f
C1723 a_2472_1562# enable 0.08694f
C1724 a_26296_2002# enable 0.05124f
C1725 a_8_1562# a_992_2122# 0.07055f
C1726 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_0.gated_control 0.23535f
C1727 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[9] 1.17576f
C1728 a_46620_1580# d_out 0
C1729 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C1730 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] 0.11433f
C1731 a_46152_1562# d_out 0
C1732 a_20056_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C1733 ShiftReg_row_10_2$1_0.Q[1] phi_1 0.05798f
C1734 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C1735 a_31208_1562# phi_1 0.70141f
C1736 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C1737 a_38776_2002# pin 0.00117f
C1738 a_24968_1562# a_27432_1562# 0
C1739 ShiftReg_row_10_2$1_0.Q[4] ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C1740 a_22176_2122# phi_2 0.04011f
C1741 a_3800_2002# swmatrix_Tgate_9.gated_control 0.01014f
C1742 a_53376_2122# enable 0.11443f
C1743 a_19712_2122# phi_2 0.04895f
C1744 a_50912_2122# enable 0.11055f
C1745 a_51116_2122# vdd 0.01506f
C1746 a_32536_2002# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1747 a_50764_1577# swmatrix_Tgate_1.gated_control 0
C1748 ShiftReg_row_10_2$1_0.Q[9] a_56168_1562# 0.16779f
C1749 a_46988_1577# BUS[8] 0
C1750 a_35000_2002# ShiftReg_row_10_2$1_0.Q[6] 0.25874f
C1751 a_31208_1562# swmatrix_Tgate_6.gated_control 0.01446f
C1752 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_34656_2122# 0.01536f
C1753 a_37448_1562# phi_2 0.02762f
C1754 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1755 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C1756 swmatrix_Tgate_8.gated_control a_12956_1580# 0
C1757 a_59616_2122# a_59820_2122# 0.01151f
C1758 a_12488_1562# a_13816_2002# 0.02403f
C1759 a_59100_1580# a_59468_2122# 0.00294f
C1760 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C1761 a_3456_2122# a_3700_1577# 0.01595f
C1762 a_58632_1562# a_57496_2002# 0
C1763 a_28760_2002# enable 0.0522f
C1764 ShiftReg_row_10_2$1_0.Q[5] vdd 0.57782f
C1765 a_57152_2122# a_57004_2122# 0
C1766 a_25436_1580# enable 0.05108f
C1767 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00721f
C1768 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C1769 a_7576_2002# vdd 0.32602f
C1770 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_22520_2002# 0.00242f
C1771 a_47136_2122# d_out 0
C1772 a_48601_1539# phi_2 0
C1773 a_19196_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0
C1774 a_992_2122# BUS[1] 0.01984f
C1775 a_47480_2002# a_47340_2122# 0.00109f
C1776 a_41240_2002# pin 0.00147f
C1777 a_44672_2122# a_44524_1577# 0
C1778 a_1196_2122# enable 0.00368f
C1779 a_44156_1580# a_44524_2122# 0.00294f
C1780 phi_1 D_in 0.02231f
C1781 a_37916_1580# pin 0
C1782 a_29881_1539# BUS[5] 0
C1783 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C1784 a_24968_1562# a_25952_2122# 0.07055f
C1785 a_53580_2122# vdd 0.01506f
C1786 a_2940_1580# swmatrix_Tgate_9.gated_control 0.00668f
C1787 swmatrix_Tgate_1.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C1788 a_50764_2122# vdd 0.00491f
C1789 swmatrix_Tgate_0.gated_control BUS[6] 0.00677f
C1790 a_35000_2002# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C1791 vdd pin 9.80638f
C1792 a_46620_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1793 a_31676_1580# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1794 a_46152_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1795 ShiftReg_row_10_2$1_0.Q[8] phi_1 0.05798f
C1796 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C1797 a_8_1562# vdd 1.0074f
C1798 a_51156_1577# swmatrix_Tgate_1.gated_control 0
C1799 a_22520_2002# d_out 0
C1800 a_51116_2122# swmatrix_Tgate_1.gated_control 0
C1801 a_34140_1580# ShiftReg_row_10_2$1_0.Q[6] 0.00101f
C1802 a_47380_1577# BUS[8] 0
C1803 a_33672_1562# ShiftReg_row_10_2$1_0.Q[6] 0.00225f
C1804 a_32536_2002# a_32436_1577# 0
C1805 a_31676_1580# a_32044_1577# 0.00194f
C1806 a_59616_2122# a_59468_2122# 0
C1807 enable BUS[2] 0.21339f
C1808 a_32536_2002# a_32396_2122# 0.00109f
C1809 a_59100_1580# a_59960_2002# 0.00888f
C1810 a_12488_1562# a_12956_1580# 0.30528f
C1811 phi_1 BUS[9] 0.09482f
C1812 a_58632_1562# a_59960_2002# 0.02403f
C1813 a_57152_2122# a_57496_2002# 0.57845f
C1814 a_58632_1562# a_56636_1580# 0
C1815 a_27900_1580# enable 0.05124f
C1816 a_27432_1562# enable 0.08694f
C1817 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00327f
C1818 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_1.gated_control 0.33472f
C1819 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C1820 a_61081_1539# phi_2 0
C1821 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_0.gated_control 0.22418f
C1822 ShiftReg_row_10_2$1_0.Q[9] phi_2 0.63578f
C1823 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_1 0.01369f
C1824 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_21660_1580# 0.36162f
C1825 a_6716_1580# vdd 0.42253f
C1826 a_46988_1577# phi_2 0
C1827 swmatrix_Tgate_4.gated_control swmatrix_Tgate_7.gated_control 0.01259f
C1828 a_6248_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C1829 swmatrix_Tgate_8.gated_control phi_2 0.31092f
C1830 swmatrix_Tgate_9.gated_control a_4921_1539# 0.00113f
C1831 a_21192_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.16689f
C1832 a_1336_2002# pin 0.00136f
C1833 a_44672_2122# a_44916_1577# 0.01595f
C1834 a_40380_1580# pin 0
C1835 swmatrix_Tgate_0.gated_control enable 0.50853f
C1836 a_44672_2122# a_44876_2122# 0.01151f
C1837 a_39912_1562# pin 0.00214f
C1838 a_44156_1580# a_45016_2002# 0.00888f
C1839 a_28268_1577# BUS[5] 0
C1840 a_8_1562# a_1336_2002# 0.02403f
C1841 a_992_2122# a_476_1580# 0.30053f
C1842 a_38284_1577# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1843 a_3456_2122# swmatrix_Tgate_9.gated_control 0.01553f
C1844 ShiftReg_row_10_2$1_0.Q[8] ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C1845 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[8] 1.17576f
C1846 a_53228_2122# vdd 0.00491f
C1847 a_34140_1580# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C1848 swmatrix_Tgate_2.gated_control BUS[10] 0.86839f
C1849 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_46988_1577# 0
C1850 a_844_2122# BUS[1] 0
C1851 a_51256_2002# vdd 0.32602f
C1852 a_47136_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C1853 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C1854 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_5.gated_control 0.23535f
C1855 a_33672_1562# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C1856 phi_1 d_out 0.10096f
C1857 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C1858 a_21660_1580# d_out 0
C1859 a_53580_2122# swmatrix_Tgate_1.gated_control 0
C1860 a_21192_1562# d_out 0
C1861 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C1862 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[9] 0.10641f
C1863 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] 0.11433f
C1864 swmatrix_Tgate_1.gated_control pin 1.20655f
C1865 a_13816_2002# pin 0.00117f
C1866 a_12488_1562# a_14952_1562# 0
C1867 a_59616_2122# a_59960_2002# 0.57845f
C1868 vdd BUS[1] 0.59166f
C1869 ShiftReg_row_10_2$1_0.Q[2] ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.08575f
C1870 a_58632_1562# a_59100_1580# 0.30528f
C1871 a_844_1577# enable 0.00235f
C1872 a_28416_2122# enable 0.11443f
C1873 a_57152_2122# a_56636_1580# 0.30053f
C1874 a_25952_2122# enable 0.11055f
C1875 a_12488_1562# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1876 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_56168_1562# 0
C1877 a_26156_2122# vdd 0.01506f
C1878 a_59468_1577# phi_2 0
C1879 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN D_in 0
C1880 swmatrix_Tgate_6.gated_control d_out 0.35904f
C1881 a_38284_1577# swmatrix_Tgate_0.gated_control 0
C1882 ShiftReg_row_10_2$1_0.Q[7] a_43688_1562# 0.16779f
C1883 a_11161_1539# BUS[2] 0
C1884 a_22520_2002# ShiftReg_row_10_2$1_0.Q[4] 0.25874f
C1885 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_8.gated_control 0.17173f
C1886 a_50764_1577# phi_2 0
C1887 a_47380_1577# phi_2 0
C1888 a_18728_1562# swmatrix_Tgate_7.gated_control 0.01446f
C1889 a_8712_1562# vdd 1.04286f
C1890 swmatrix_Tgate_9.gated_control a_3308_1577# 0
C1891 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_22176_2122# 0.01536f
C1892 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.43061f
C1893 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1894 swmatrix_Tgate_7.gated_control BUS[3] 0.00677f
C1895 a_12488_1562# phi_2 0.02762f
C1896 a_47136_2122# a_47340_2122# 0.01151f
C1897 a_46620_1580# a_46988_2122# 0.00294f
C1898 a_40896_2122# pin 0.00304f
C1899 a_43688_1562# enable 0.08752f
C1900 a_46152_1562# a_45016_2002# 0
C1901 a_38676_1577# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1902 a_992_2122# a_2472_1562# 0.00268f
C1903 a_38432_2122# pin 0
C1904 a_44672_2122# a_44524_2122# 0
C1905 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C1906 a_28660_1577# BUS[5] 0
C1907 ShiftReg_row_10_2$1_0.Q[8] a_48601_1539# 0.00241f
C1908 a_53720_2002# vdd 0.3289f
C1909 a_34656_2122# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C1910 a_32192_2122# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1911 a_50396_1580# vdd 0.42253f
C1912 a_1336_2002# BUS[1] 0.01222f
C1913 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_10040_2002# 0.00242f
C1914 a_22176_2122# d_out 0
C1915 a_23641_1539# phi_2 0
C1916 a_56168_1562# pin 0.00162f
C1917 a_51256_2002# swmatrix_Tgate_1.gated_control 0.01141f
C1918 a_476_1580# a_844_2122# 0.00294f
C1919 a_35000_2002# a_34860_2122# 0.00109f
C1920 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.09501f
C1921 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1922 a_54841_1539# enable 0.00398f
C1923 a_44876_2122# phi_1 0.00534f
C1924 pin BUS[8] 10.5929f
C1925 a_16280_2002# pin 0.00147f
C1926 a_32192_2122# a_32044_1577# 0
C1927 a_31676_1580# a_32044_2122# 0.00294f
C1928 a_12956_1580# pin 0
C1929 a_12488_1562# a_13472_2122# 0.07055f
C1930 a_59616_2122# a_59100_1580# 0.30053f
C1931 a_1236_1577# enable 0.00582f
C1932 a_58632_1562# a_59616_2122# 0.07055f
C1933 a_57152_2122# a_58632_1562# 0.00268f
C1934 a_28620_2122# vdd 0.01506f
C1935 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C1936 a_25804_2122# vdd 0.00491f
C1937 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C1938 a_59860_1577# phi_2 0
C1939 a_34140_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1940 a_476_1580# vdd 0.42253f
C1941 ShiftReg_row_10_2$1_0.Q[4] phi_1 0.05798f
C1942 a_9548_1577# BUS[2] 0
C1943 a_33672_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C1944 a_38676_1577# swmatrix_Tgate_0.gated_control 0
C1945 a_7232_2122# vdd 0.56061f
C1946 swmatrix_Tgate_9.gated_control a_7084_1577# 0
C1947 a_21660_1580# ShiftReg_row_10_2$1_0.Q[4] 0.00101f
C1948 a_38636_2122# swmatrix_Tgate_0.gated_control 0
C1949 a_51156_1577# phi_2 0
C1950 a_20056_2002# a_19956_1577# 0
C1951 a_21192_1562# ShiftReg_row_10_2$1_0.Q[4] 0.00225f
C1952 a_19196_1580# a_19564_1577# 0.00194f
C1953 swmatrix_Tgate_9.gated_control a_3700_1577# 0
C1954 a_51116_2122# phi_2 0.00411f
C1955 a_46620_1580# a_47480_2002# 0.00888f
C1956 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1957 a_47136_2122# a_46988_2122# 0
C1958 a_20056_2002# a_19916_2122# 0.00109f
C1959 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C1960 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C1961 a_46152_1562# a_47480_2002# 0.02403f
C1962 a_46152_1562# a_44156_1580# 0
C1963 a_44672_2122# a_45016_2002# 0.57845f
C1964 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[6] 0.10641f
C1965 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_0.gated_control 0.33472f
C1966 a_48601_1539# d_out 0
C1967 a_52860_1580# vdd 0.4252f
C1968 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C1969 a_52392_1562# vdd 1.04286f
C1970 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_5.gated_control 0.22418f
C1971 ShiftReg_row_10_2$1_0.Q[5] phi_2 0.63578f
C1972 a_22028_1577# phi_2 0
C1973 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_9180_1580# 0.36162f
C1974 ShiftReg_row_10_2$1_0.Q[9] BUS[9] 0.0247f
C1975 a_47340_2122# phi_1 0.00477f
C1976 a_53720_2002# swmatrix_Tgate_1.gated_control 0.01014f
C1977 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C1978 a_44524_2122# phi_1 0.00201f
C1979 a_53228_1577# enable 0.0022f
C1980 a_992_2122# a_1196_2122# 0.01151f
C1981 a_476_1580# a_1336_2002# 0.00888f
C1982 a_50396_1580# swmatrix_Tgate_1.gated_control 0.00829f
C1983 a_15420_1580# pin 0
C1984 a_32192_2122# a_32436_1577# 0.01595f
C1985 swmatrix_Tgate_4.gated_control enable 0.50853f
C1986 a_31676_1580# a_32536_2002# 0.00888f
C1987 a_14952_1562# pin 0.00214f
C1988 a_32192_2122# a_32396_2122# 0.01151f
C1989 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C1990 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[7] 1.17576f
C1991 a_3660_2122# enable 0.00368f
C1992 a_7576_2002# phi_2 0.03207f
C1993 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C1994 ShiftReg_row_10_2$1_0.Q[6] ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C1995 a_28268_2122# vdd 0.00491f
C1996 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_34508_1577# 0
C1997 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_4.gated_control 0.23535f
C1998 a_2472_1562# vdd 1.04253f
C1999 a_26296_2002# vdd 0.32602f
C2000 swmatrix_Tgate_2.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00605f
C2001 a_34656_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C2002 a_9940_1577# BUS[2] 0
C2003 a_41100_2122# swmatrix_Tgate_0.gated_control 0
C2004 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] 0.11433f
C2005 swmatrix_Tgate_5.gated_control pin 1.20655f
C2006 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C2007 a_53580_2122# phi_2 0.00422f
C2008 phi_2 pin 0.18641f
C2009 a_50764_2122# phi_2 0
C2010 a_47136_2122# a_47480_2002# 0.57845f
C2011 a_61081_1539# d_out 0.00256f
C2012 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34484f
C2013 a_46152_1562# a_46620_1580# 0.30528f
C2014 a_44672_2122# a_44156_1580# 0.30053f
C2015 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C2016 a_8_1562# phi_2 0.03129f
C2017 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_43688_1562# 0
C2018 ShiftReg_row_10_2$1_0.Q[9] d_out 0
C2019 a_38776_2002# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2020 a_46988_1577# d_out 0
C2021 ShiftReg_row_10_2$1_0.Q[8] a_50764_1577# 0
C2022 swmatrix_Tgate_8.gated_control d_out 0.35904f
C2023 a_53376_2122# vdd 0.56003f
C2024 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C2025 swmatrix_Tgate_0.gated_control BUS[7] 0.86839f
C2026 ShiftReg_row_10_2$1_0.Q[5] a_31208_1562# 0.16779f
C2027 a_50912_2122# vdd 0.56061f
C2028 a_25804_1577# swmatrix_Tgate_5.gated_control 0
C2029 a_10040_2002# ShiftReg_row_10_2$1_0.Q[2] 0.25874f
C2030 a_25804_1577# phi_2 0
C2031 a_46988_2122# phi_1 0.00164f
C2032 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_9696_2122# 0.01536f
C2033 a_22420_1577# phi_2 0
C2034 a_45016_2002# phi_1 0.01314f
C2035 a_52860_1580# swmatrix_Tgate_1.gated_control 0.00668f
C2036 a_57004_1577# enable 0.0022f
C2037 a_34140_1580# a_34508_2122# 0.00294f
C2038 a_53620_1577# enable 0.00579f
C2039 a_34656_2122# a_34860_2122# 0.01151f
C2040 a_52392_1562# swmatrix_Tgate_1.gated_control 0.00985f
C2041 a_2472_1562# a_1336_2002# 0
C2042 a_18728_1562# enable 0.08752f
C2043 a_15936_2122# pin 0.00304f
C2044 ShiftReg_row_10_2$1_0.Q[1] a_7576_2002# 0.00242f
C2045 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_48601_1539# 0.0097f
C2046 a_33672_1562# a_32536_2002# 0
C2047 a_13472_2122# pin 0
C2048 a_6716_1580# phi_2 0.03321f
C2049 a_32192_2122# a_32044_2122# 0
C2050 enable BUS[3] 0.21339f
C2051 a_3308_2122# enable 0.00101f
C2052 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D d_out 0
C2053 phi_1 BUS[10] 0.09482f
C2054 ShiftReg_row_10_2$1_0.Q[6] a_36121_1539# 0.00241f
C2055 a_28760_2002# vdd 0.3289f
C2056 a_1336_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.2556f
C2057 a_25436_1580# vdd 0.42253f
C2058 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D BUS[3] 0.10641f
C2059 ShiftReg_row_10_2$1_0.Q[1] pin 0.01551f
C2060 a_38776_2002# swmatrix_Tgate_0.gated_control 0.01141f
C2061 a_53228_2122# phi_2 0
C2062 a_22520_2002# a_22380_2122# 0.00109f
C2063 a_31208_1562# pin 0.00162f
C2064 a_19916_2122# phi_1 0.00534f
C2065 a_29881_1539# enable 0.00398f
C2066 a_51256_2002# phi_2 0.03207f
C2067 a_19712_2122# a_19564_1577# 0
C2068 a_19196_1580# a_19564_2122# 0.00294f
C2069 a_47136_2122# a_46620_1580# 0.30053f
C2070 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00355f
C2071 a_59468_1577# d_out 0
C2072 a_844_1577# a_992_2122# 0
C2073 a_46152_1562# a_47136_2122# 0.07055f
C2074 ShiftReg_row_10_2$1_0.Q[6] BUS[6] 0.0247f
C2075 a_1196_2122# vdd 0.01506f
C2076 a_44672_2122# a_46152_1562# 0.00268f
C2077 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_1 0.02073f
C2078 a_41240_2002# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00155f
C2079 a_37916_1580# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2080 a_21660_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C2081 a_47380_1577# d_out 0
C2082 phi_2 BUS[1] 0.10922f
C2083 a_21192_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C2084 a_26196_1577# swmatrix_Tgate_5.gated_control 0
C2085 a_26156_2122# swmatrix_Tgate_5.gated_control 0
C2086 a_9180_1580# ShiftReg_row_10_2$1_0.Q[2] 0.00101f
C2087 a_26196_1577# phi_2 0
C2088 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vdd 4.98668f
C2089 a_26156_2122# phi_2 0.00411f
C2090 a_47480_2002# phi_1 0.01261f
C2091 a_51156_1577# BUS[9] 0
C2092 a_53376_2122# swmatrix_Tgate_1.gated_control 0.01553f
C2093 a_57396_1577# enable 0.00577f
C2094 a_57356_2122# enable 0.00368f
C2095 a_34656_2122# a_34508_2122# 0
C2096 a_34140_1580# a_35000_2002# 0.00888f
C2097 a_50912_2122# swmatrix_Tgate_1.gated_control 0.01538f
C2098 a_51116_2122# BUS[9] 0
C2099 a_44156_1580# phi_1 0.0533f
C2100 a_33672_1562# a_35000_2002# 0.02403f
C2101 a_6248_1562# swmatrix_Tgate_9.gated_control 0.00493f
C2102 ShiftReg_row_10_2$1_0.Q[1] a_6716_1580# 0.36203f
C2103 swmatrix_Tgate_2.gated_control phi_1 0.00906f
C2104 a_32192_2122# a_32536_2002# 0.57845f
C2105 a_33672_1562# a_31676_1580# 0
C2106 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_5.gated_control 0.33472f
C2107 vdd BUS[2] 0.58892f
C2108 a_8712_1562# phi_2 0.60119f
C2109 a_3800_2002# enable 0.0522f
C2110 a_23641_1539# d_out 0
C2111 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I phi_2 0.03773f
C2112 a_27900_1580# vdd 0.4252f
C2113 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_4.gated_control 0.22418f
C2114 a_27432_1562# vdd 1.04286f
C2115 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[9] 0
C2116 a_1336_2002# a_1196_2122# 0.00109f
C2117 ShiftReg_row_10_2$1_0.Q[6] enable 0.513f
C2118 a_41240_2002# swmatrix_Tgate_0.gated_control 0.01014f
C2119 a_22380_2122# phi_1 0.00477f
C2120 a_19564_2122# phi_1 0.00201f
C2121 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[6] 1.17576f
C2122 a_37916_1580# swmatrix_Tgate_0.gated_control 0.00829f
C2123 a_53720_2002# phi_2 0.03174f
C2124 a_28268_1577# enable 0.0022f
C2125 a_50396_1580# phi_2 0.03321f
C2126 swmatrix_Tgate_7.gated_control BUS[4] 0.86839f
C2127 D_in pin 0.00658f
C2128 a_19712_2122# a_19956_1577# 0.01595f
C2129 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN d_out 0.46167f
C2130 a_19712_2122# a_19916_2122# 0.01151f
C2131 a_19196_1580# a_20056_2002# 0.00888f
C2132 a_44524_1577# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2133 a_59860_1577# d_out 0
C2134 a_7084_2122# enable 0.00101f
C2135 a_1236_1577# a_992_2122# 0.01595f
C2136 ShiftReg_row_10_2$1_0.Q[4] ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C2137 swmatrix_Tgate_0.gated_control vdd 1.8044f
C2138 a_8_1562# D_in 0.15891f
C2139 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_22028_1577# 0
C2140 a_40380_1580# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00173f
C2141 a_22176_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C2142 ShiftReg_row_10_2$1_0.Q[1] BUS[1] 0.01648f
C2143 a_39912_1562# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.0046f
C2144 ShiftReg_row_10_2$1_0.Q[8] pin 0.01625f
C2145 a_28620_2122# swmatrix_Tgate_5.gated_control 0
C2146 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D enable 0.20415f
C2147 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] 0.11433f
C2148 a_28620_2122# phi_2 0.00422f
C2149 a_476_1580# phi_2 0.03488f
C2150 a_59820_2122# enable 0.00368f
C2151 a_46620_1580# phi_1 0.01277f
C2152 a_53580_2122# BUS[9] 0.00104f
C2153 a_25804_2122# phi_2 0
C2154 a_57004_2122# enable 0.00101f
C2155 a_46152_1562# phi_1 0.01733f
C2156 pin BUS[9] 10.5929f
C2157 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C2158 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C2159 a_34656_2122# a_35000_2002# 0.57845f
C2160 a_33672_1562# a_34140_1580# 0.30528f
C2161 a_18728_1562# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2162 a_32192_2122# a_31676_1580# 0.30053f
C2163 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN pin 1.45295f
C2164 a_7232_2122# phi_2 0.04895f
C2165 ShiftReg_row_10_2$1_0.Q[5] d_out 0
C2166 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_31208_1562# 0
C2167 a_2940_1580# enable 0.05124f
C2168 ShiftReg_row_10_2$1_0.Q[6] a_38284_1577# 0
C2169 a_22028_1577# d_out 0
C2170 a_28416_2122# vdd 0.56003f
C2171 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN enable 0.09895f
C2172 a_25952_2122# vdd 0.56061f
C2173 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D pin 0.00147f
C2174 a_13324_1577# swmatrix_Tgate_4.gated_control 0
C2175 ShiftReg_row_10_2$1_0.Q[3] a_18728_1562# 0.16779f
C2176 ShiftReg_row_10_2$1_0.Q[3] BUS[3] 0.0247f
C2177 a_22028_2122# phi_1 0.00164f
C2178 a_40380_1580# swmatrix_Tgate_0.gated_control 0.00668f
C2179 a_22176_2122# a_22380_2122# 0.01151f
C2180 a_32044_1577# enable 0.0022f
C2181 a_20056_2002# phi_1 0.01314f
C2182 a_21660_1580# a_22028_2122# 0.00294f
C2183 a_39912_1562# swmatrix_Tgate_0.gated_control 0.00985f
C2184 a_28660_1577# enable 0.00579f
C2185 a_52860_1580# phi_2 0.07395f
C2186 a_52392_1562# phi_2 0.60119f
C2187 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_36121_1539# 0.0097f
C2188 a_21192_1562# a_20056_2002# 0
C2189 a_19712_2122# a_19564_2122# 0
C2190 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.90801f
C2191 a_44916_1577# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2192 a_32436_1577# BUS[6] 0
C2193 a_43688_1562# vdd 1.00072f
C2194 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_1 0
C2195 ShiftReg_row_10_2$1_0.Q[4] a_23641_1539# 0.00241f
C2196 a_40896_2122# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00387f
C2197 a_32396_2122# BUS[6] 0
C2198 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C2199 d_out pin 1.8694f
C2200 a_38432_2122# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2201 a_44524_1577# pin 0
C2202 a_61081_1539# BUS[10] 0
C2203 ShiftReg_row_10_2$1_0.Q[8] a_51256_2002# 0.00242f
C2204 D_in BUS[1] 0
C2205 a_41140_1577# pin 0
C2206 a_28268_2122# phi_2 0
C2207 a_4921_1539# enable 0.00398f
C2208 a_26296_2002# swmatrix_Tgate_5.gated_control 0.01141f
C2209 a_10040_2002# a_9900_2122# 0.00109f
C2210 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2211 a_26296_2002# phi_2 0.03207f
C2212 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[6] 0
C2213 a_53228_2122# BUS[9] 0
C2214 a_47136_2122# phi_1 0.01804f
C2215 a_59468_2122# enable 0.00101f
C2216 a_2472_1562# phi_2 0.60119f
C2217 a_34656_2122# a_34140_1580# 0.30053f
C2218 a_51256_2002# BUS[9] 0.01182f
C2219 a_44672_2122# phi_1 0.01882f
C2220 a_57496_2002# enable 0.05124f
C2221 ShiftReg_row_10_2$1_0.Q[1] a_7232_2122# 0.01552f
C2222 a_33672_1562# a_34656_2122# 0.07055f
C2223 a_32192_2122# a_33672_1562# 0.00268f
C2224 a_3456_2122# enable 0.11443f
C2225 a_22420_1577# d_out 0
C2226 a_9180_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0
C2227 a_13716_1577# swmatrix_Tgate_4.gated_control 0
C2228 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D phi_2 0.45413f
C2229 a_13676_2122# swmatrix_Tgate_4.gated_control 0
C2230 a_32436_1577# enable 0.00577f
C2231 a_22520_2002# phi_1 0.01261f
C2232 a_40896_2122# swmatrix_Tgate_0.gated_control 0.01553f
C2233 a_22176_2122# a_22028_2122# 0
C2234 a_32396_2122# enable 0.00368f
C2235 a_21660_1580# a_22520_2002# 0.00888f
C2236 a_19196_1580# phi_1 0.0533f
C2237 a_38432_2122# swmatrix_Tgate_0.gated_control 0.01538f
C2238 a_53376_2122# phi_2 0.04011f
C2239 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.00126f
C2240 a_21192_1562# a_22520_2002# 0.02403f
C2241 a_19712_2122# a_20056_2002# 0.57845f
C2242 a_21192_1562# a_19196_1580# 0
C2243 a_50912_2122# phi_2 0.04895f
C2244 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I swmatrix_Tgate_4.gated_control 0.33472f
C2245 a_34860_2122# BUS[6] 0.00104f
C2246 swmatrix_Tgate_2.gated_control a_61081_1539# 0.00113f
C2247 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I enable 0.65271f
C2248 a_59468_1577# BUS[10] 0
C2249 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_2.gated_control 0.17173f
C2250 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN BUS[5] 1.17576f
C2251 a_49928_1562# swmatrix_Tgate_3.gated_control 0.00493f
C2252 ShiftReg_row_10_2$1_0.Q[8] a_50396_1580# 0.36203f
C2253 ShiftReg_row_10_2$1_0.Q[2] enable 0.513f
C2254 a_28760_2002# swmatrix_Tgate_5.gated_control 0.01014f
C2255 a_28760_2002# phi_2 0.03174f
C2256 a_25436_1580# swmatrix_Tgate_5.gated_control 0.00829f
C2257 a_1236_1577# a_1336_2002# 0
C2258 a_3308_1577# enable 0.0022f
C2259 ShiftReg_row_10_2$1_0.Q[1] a_2472_1562# 0.00225f
C2260 a_476_1580# D_in 0.36155f
C2261 a_25436_1580# phi_2 0.03321f
C2262 a_59960_2002# enable 0.0522f
C2263 a_53720_2002# BUS[9] 0.00972f
C2264 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vdd 0.42786f
C2265 a_50396_1580# BUS[9] 0.0049f
C2266 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[1] 0
C2267 a_56636_1580# enable 0.05108f
C2268 d_out BUS[1] 0.16227f
C2269 swmatrix_Tgate_4.gated_control vdd 1.8044f
C2270 enable BUS[4] 0.21339f
C2271 ShiftReg_row_10_2$1_0.Q[2] ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01068f
C2272 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I pin 0
C2273 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D a_9548_1577# 0
C2274 a_3660_2122# vdd 0.01506f
C2275 ShiftReg_row_10_2$1_0.Q[1] ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.01102f
C2276 swmatrix_Tgate_1.gated_control a_54841_1539# 0.00113f
C2277 a_56168_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D 0.00116f
C2278 a_9696_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I 0.00144f
C2279 ShiftReg_row_10_2$1_0.Q[4] pin 0.01625f
C2280 a_16140_2122# swmatrix_Tgate_4.gated_control 0
C2281 a_1196_2122# phi_2 0.00411f
C2282 a_13716_1577# BUS[3] 0
C2283 a_13676_2122# BUS[3] 0
C2284 a_8712_1562# d_out 0
C2285 a_34860_2122# enable 0.00368f
C2286 a_21660_1580# phi_1 0.01277f
C2287 a_32044_2122# enable 0.00101f
C2288 a_22176_2122# a_22520_2002# 0.57845f
C2289 a_21192_1562# phi_1 0.01733f
C2290 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I d_out 0
C2291 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vdd 0.34531f
C2292 a_21192_1562# a_21660_1580# 0.30528f
C2293 a_19712_2122# a_19196_1580# 0.30053f
C2294 a_45016_2002# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0
C2295 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I a_18728_1562# 0
C2296 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN phi_2 0.00159f
C2297 ShiftReg_row_10_2$1_0.Q[4] a_25804_1577# 0
C2298 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I BUS[3] 0
C2299 a_34508_2122# BUS[6] 0
C2300 BUS[10] vss 3.81451f
C2301 BUS[9] vss 3.81467f
C2302 BUS[8] vss 3.81467f
C2303 BUS[7] vss 3.81467f
C2304 BUS[6] vss 3.81467f
C2305 BUS[5] vss 3.81467f
C2306 BUS[4] vss 3.81467f
C2307 BUS[3] vss 3.81467f
C2308 BUS[2] vss 3.81467f
C2309 BUS[1] vss 3.81197f
C2310 pin vss 24.20904f
C2311 d_out vss 32.05165f
C2312 enable vss 24.5348f
C2313 phi_2 vss 21.36711f
C2314 D_in vss 0.46366f
C2315 phi_1 vss 31.70718f
C2316 vdd vss 0.30382p
C2317 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.68096f
C2318 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2319 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2320 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2321 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2322 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2323 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2324 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.6793f
C2325 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.67985f
C2326 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN vss 1.67536f
C2327 a_61081_1539# vss 0.0072f
C2328 a_59468_1577# vss 0.0042f
C2329 a_59860_1577# vss 0.0095f
C2330 swmatrix_Tgate_2.gated_control vss 3.0993f
C2331 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.77346f
C2332 a_57004_1577# vss 0.0042f
C2333 a_57396_1577# vss 0.0095f
C2334 a_59960_2002# vss 0.4183f
C2335 a_59100_1580# vss 0.52809f
C2336 a_59616_2122# vss 1.12791f
C2337 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2338 a_54841_1539# vss 0.0072f
C2339 a_53228_1577# vss 0.0042f
C2340 a_53620_1577# vss 0.0095f
C2341 a_57496_2002# vss 0.42106f
C2342 a_56636_1580# vss 0.53029f
C2343 a_58632_1562# vss 1.18034f
C2344 a_57152_2122# vss 1.14755f
C2345 swmatrix_Tgate_1.gated_control vss 3.08335f
C2346 a_56168_1562# vss 1.18379f
C2347 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2348 ShiftReg_row_10_2$1_0.Q[9] vss 1.42244f
C2349 a_50764_1577# vss 0.0042f
C2350 a_51156_1577# vss 0.0095f
C2351 a_53720_2002# vss 0.4183f
C2352 a_52860_1580# vss 0.52809f
C2353 a_53376_2122# vss 1.12791f
C2354 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2355 a_48601_1539# vss 0.0072f
C2356 a_46988_1577# vss 0.0042f
C2357 a_47380_1577# vss 0.0095f
C2358 a_51256_2002# vss 0.42106f
C2359 a_50396_1580# vss 0.53029f
C2360 a_52392_1562# vss 1.18034f
C2361 a_50912_2122# vss 1.14755f
C2362 swmatrix_Tgate_3.gated_control vss 3.08335f
C2363 a_49928_1562# vss 1.18379f
C2364 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2365 ShiftReg_row_10_2$1_0.Q[8] vss 1.42244f
C2366 a_44524_1577# vss 0.0042f
C2367 a_44916_1577# vss 0.0095f
C2368 a_47480_2002# vss 0.4183f
C2369 a_46620_1580# vss 0.52809f
C2370 a_47136_2122# vss 1.12791f
C2371 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2372 a_42361_1539# vss 0.0072f
C2373 a_40748_1577# vss 0.0042f
C2374 a_41140_1577# vss 0.0095f
C2375 a_45016_2002# vss 0.42106f
C2376 a_44156_1580# vss 0.53029f
C2377 a_46152_1562# vss 1.18034f
C2378 a_44672_2122# vss 1.14755f
C2379 swmatrix_Tgate_0.gated_control vss 3.08335f
C2380 a_43688_1562# vss 1.18379f
C2381 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2382 ShiftReg_row_10_2$1_0.Q[7] vss 1.42244f
C2383 a_38284_1577# vss 0.0042f
C2384 a_38676_1577# vss 0.0095f
C2385 a_41240_2002# vss 0.4183f
C2386 a_40380_1580# vss 0.52809f
C2387 a_40896_2122# vss 1.12791f
C2388 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2389 a_36121_1539# vss 0.0072f
C2390 a_34508_1577# vss 0.0042f
C2391 a_34900_1577# vss 0.0095f
C2392 a_38776_2002# vss 0.42106f
C2393 a_37916_1580# vss 0.53029f
C2394 a_39912_1562# vss 1.18034f
C2395 a_38432_2122# vss 1.14755f
C2396 swmatrix_Tgate_6.gated_control vss 3.08335f
C2397 a_37448_1562# vss 1.18379f
C2398 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2399 ShiftReg_row_10_2$1_0.Q[6] vss 1.42244f
C2400 a_32044_1577# vss 0.0042f
C2401 a_32436_1577# vss 0.0095f
C2402 a_35000_2002# vss 0.4183f
C2403 a_34140_1580# vss 0.52809f
C2404 a_34656_2122# vss 1.12791f
C2405 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2406 a_29881_1539# vss 0.0072f
C2407 a_28268_1577# vss 0.0042f
C2408 a_28660_1577# vss 0.0095f
C2409 a_32536_2002# vss 0.42106f
C2410 a_31676_1580# vss 0.53029f
C2411 a_33672_1562# vss 1.18034f
C2412 a_32192_2122# vss 1.14755f
C2413 swmatrix_Tgate_5.gated_control vss 3.08335f
C2414 a_31208_1562# vss 1.18379f
C2415 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2416 ShiftReg_row_10_2$1_0.Q[5] vss 1.42244f
C2417 a_25804_1577# vss 0.0042f
C2418 a_26196_1577# vss 0.0095f
C2419 a_28760_2002# vss 0.4183f
C2420 a_27900_1580# vss 0.52809f
C2421 a_28416_2122# vss 1.12791f
C2422 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2423 a_23641_1539# vss 0.0072f
C2424 a_22028_1577# vss 0.0042f
C2425 a_22420_1577# vss 0.0095f
C2426 a_26296_2002# vss 0.42106f
C2427 a_25436_1580# vss 0.53029f
C2428 a_27432_1562# vss 1.18034f
C2429 a_25952_2122# vss 1.14755f
C2430 swmatrix_Tgate_7.gated_control vss 3.08335f
C2431 a_24968_1562# vss 1.18379f
C2432 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2433 ShiftReg_row_10_2$1_0.Q[4] vss 1.42244f
C2434 a_19564_1577# vss 0.0042f
C2435 a_19956_1577# vss 0.0095f
C2436 a_22520_2002# vss 0.4183f
C2437 a_21660_1580# vss 0.52809f
C2438 a_22176_2122# vss 1.12791f
C2439 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2440 a_17401_1539# vss 0.0072f
C2441 a_15788_1577# vss 0.0042f
C2442 a_16180_1577# vss 0.0095f
C2443 a_20056_2002# vss 0.42106f
C2444 a_19196_1580# vss 0.53029f
C2445 a_21192_1562# vss 1.18034f
C2446 a_19712_2122# vss 1.14755f
C2447 swmatrix_Tgate_4.gated_control vss 3.08335f
C2448 a_18728_1562# vss 1.18379f
C2449 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2450 ShiftReg_row_10_2$1_0.Q[3] vss 1.42244f
C2451 a_13324_1577# vss 0.0042f
C2452 a_13716_1577# vss 0.0095f
C2453 a_16280_2002# vss 0.4183f
C2454 a_15420_1580# vss 0.52809f
C2455 a_15936_2122# vss 1.12791f
C2456 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2457 a_11161_1539# vss 0.0072f
C2458 a_9548_1577# vss 0.0042f
C2459 a_9940_1577# vss 0.0095f
C2460 a_13816_2002# vss 0.42106f
C2461 a_12956_1580# vss 0.53029f
C2462 a_14952_1562# vss 1.18034f
C2463 a_13472_2122# vss 1.14755f
C2464 swmatrix_Tgate_8.gated_control vss 3.09123f
C2465 a_12488_1562# vss 1.18379f
C2466 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76709f
C2467 ShiftReg_row_10_2$1_0.Q[2] vss 1.42244f
C2468 a_7084_1577# vss 0.0042f
C2469 a_7476_1577# vss 0.0095f
C2470 a_10040_2002# vss 0.4183f
C2471 a_9180_1580# vss 0.52809f
C2472 a_9696_2122# vss 1.12791f
C2473 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66698f
C2474 a_4921_1539# vss 0.0072f
C2475 a_3308_1577# vss 0.0042f
C2476 a_3700_1577# vss 0.0095f
C2477 a_7576_2002# vss 0.42106f
C2478 a_6716_1580# vss 0.53029f
C2479 a_8712_1562# vss 1.18034f
C2480 a_7232_2122# vss 1.14755f
C2481 swmatrix_Tgate_9.gated_control vss 3.0913f
C2482 a_6248_1562# vss 1.18379f
C2483 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.I vss 0.76938f
C2484 ShiftReg_row_10_2$1_0.Q[1] vss 1.43147f
C2485 a_844_1577# vss 0.0042f
C2486 a_1236_1577# vss 0.0095f
C2487 a_3800_2002# vss 0.4183f
C2488 a_2940_1580# vss 0.52805f
C2489 a_3456_2122# vss 1.12761f
C2490 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1_0.D vss 0.66677f
C2491 a_1336_2002# vss 0.42099f
C2492 a_476_1580# vss 0.53043f
C2493 a_2472_1562# vss 1.18052f
C2494 a_992_2122# vss 1.14718f
C2495 a_8_1562# vss 1.18952f
C2496 d_out.t3 vss 0.06891f
C2497 d_out.t2 vss 0.08866f
C2498 d_out.n0 vss 0.08065f
C2499 d_out.n1 vss 0.04952f
C2500 d_out.n2 vss 0.20168f
C2501 d_out.t1 vss 0.08199f
C2502 d_out.t0 vss 0.05742f
C2503 d_out.n3 vss 0.09782f
C2504 BUS[7].t20 vss 0.08272f
C2505 BUS[7].t22 vss 0.08272f
C2506 BUS[7].n0 vss 0.44552f
C2507 BUS[7].t21 vss 0.08272f
C2508 BUS[7].t17 vss 0.08272f
C2509 BUS[7].n1 vss 0.44289f
C2510 BUS[7].n2 vss 0.25937f
C2511 BUS[7].t18 vss 0.08272f
C2512 BUS[7].t19 vss 0.08272f
C2513 BUS[7].n3 vss 0.44289f
C2514 BUS[7].n4 vss 0.21881f
C2515 BUS[7].t6 vss 0.66732f
C2516 BUS[7].n5 vss 0.21139f
C2517 BUS[7].t15 vss 0.08272f
C2518 BUS[7].t16 vss 0.08272f
C2519 BUS[7].n6 vss 0.44813f
C2520 BUS[7].t7 vss 0.08272f
C2521 BUS[7].t10 vss 0.08272f
C2522 BUS[7].n7 vss 0.44556f
C2523 BUS[7].n8 vss 0.25349f
C2524 BUS[7].t13 vss 0.08272f
C2525 BUS[7].t2 vss 0.08272f
C2526 BUS[7].n9 vss 0.44556f
C2527 BUS[7].n10 vss 0.14712f
C2528 BUS[7].t4 vss 0.08272f
C2529 BUS[7].t14 vss 0.08272f
C2530 BUS[7].n11 vss 0.44556f
C2531 BUS[7].n12 vss 0.14712f
C2532 BUS[7].t3 vss 0.08272f
C2533 BUS[7].t5 vss 0.08272f
C2534 BUS[7].n13 vss 0.44556f
C2535 BUS[7].n14 vss 0.14712f
C2536 BUS[7].t8 vss 0.08272f
C2537 BUS[7].t11 vss 0.08272f
C2538 BUS[7].n15 vss 0.44556f
C2539 BUS[7].n16 vss 0.14712f
C2540 BUS[7].t0 vss 0.08272f
C2541 BUS[7].t9 vss 0.08272f
C2542 BUS[7].n17 vss 0.44556f
C2543 BUS[7].n18 vss 0.14712f
C2544 BUS[7].t12 vss 0.08272f
C2545 BUS[7].t1 vss 0.08272f
C2546 BUS[7].n19 vss 0.44556f
C2547 BUS[7].n20 vss 0.11197f
C2548 BUS[7].n21 vss 0.37951f
C2549 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C2550 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C2551 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.12443f
C2552 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C2553 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C2554 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C2555 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C2556 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C2557 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C2558 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C2559 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C2560 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C2561 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C2562 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C2563 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C2564 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C2565 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C2566 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C2567 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C2568 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C2569 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C2570 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C2571 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C2572 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C2573 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C2574 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C2575 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C2576 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C2577 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C2578 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C2579 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C2580 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C2581 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C2582 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C2583 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C2584 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C2585 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C2586 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C2587 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.12443f
C2588 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C2589 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C2590 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C2591 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C2592 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C2593 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C2594 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C2595 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C2596 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C2597 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C2598 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C2599 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C2600 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C2601 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C2602 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C2603 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C2604 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C2605 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C2606 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C2607 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C2608 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C2609 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C2610 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C2611 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C2612 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C2613 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C2614 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C2615 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C2616 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C2617 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C2618 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C2619 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C2620 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C2621 BUS[9].t21 vss 0.08272f
C2622 BUS[9].t16 vss 0.08272f
C2623 BUS[9].n0 vss 0.44552f
C2624 BUS[9].t18 vss 0.08272f
C2625 BUS[9].t20 vss 0.08272f
C2626 BUS[9].n1 vss 0.44289f
C2627 BUS[9].n2 vss 0.25937f
C2628 BUS[9].t19 vss 0.08272f
C2629 BUS[9].t17 vss 0.08272f
C2630 BUS[9].n3 vss 0.44289f
C2631 BUS[9].n4 vss 0.21881f
C2632 BUS[9].t7 vss 0.66732f
C2633 BUS[9].n5 vss 0.21139f
C2634 BUS[9].t12 vss 0.08272f
C2635 BUS[9].t0 vss 0.08272f
C2636 BUS[9].n6 vss 0.44813f
C2637 BUS[9].t4 vss 0.08272f
C2638 BUS[9].t11 vss 0.08272f
C2639 BUS[9].n7 vss 0.44556f
C2640 BUS[9].n8 vss 0.25349f
C2641 BUS[9].t3 vss 0.08272f
C2642 BUS[9].t8 vss 0.08272f
C2643 BUS[9].n9 vss 0.44556f
C2644 BUS[9].n10 vss 0.14712f
C2645 BUS[9].t6 vss 0.08272f
C2646 BUS[9].t10 vss 0.08272f
C2647 BUS[9].n11 vss 0.44556f
C2648 BUS[9].n12 vss 0.14712f
C2649 BUS[9].t14 vss 0.08272f
C2650 BUS[9].t22 vss 0.08272f
C2651 BUS[9].n13 vss 0.44556f
C2652 BUS[9].n14 vss 0.14712f
C2653 BUS[9].t9 vss 0.08272f
C2654 BUS[9].t1 vss 0.08272f
C2655 BUS[9].n15 vss 0.44556f
C2656 BUS[9].n16 vss 0.14712f
C2657 BUS[9].t5 vss 0.08272f
C2658 BUS[9].t2 vss 0.08272f
C2659 BUS[9].n17 vss 0.44556f
C2660 BUS[9].n18 vss 0.14712f
C2661 BUS[9].t13 vss 0.08272f
C2662 BUS[9].t15 vss 0.08272f
C2663 BUS[9].n19 vss 0.44556f
C2664 BUS[9].n20 vss 0.11197f
C2665 BUS[9].n21 vss 0.37951f
C2666 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C2667 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C2668 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.12443f
C2669 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C2670 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C2671 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C2672 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C2673 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C2674 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C2675 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C2676 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C2677 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C2678 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C2679 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C2680 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C2681 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C2682 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C2683 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C2684 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C2685 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C2686 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C2687 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C2688 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C2689 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C2690 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C2691 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C2692 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C2693 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C2694 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C2695 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C2696 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C2697 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C2698 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C2699 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C2700 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C2701 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C2702 BUS[4].t18 vss 0.08272f
C2703 BUS[4].t19 vss 0.08272f
C2704 BUS[4].n0 vss 0.44552f
C2705 BUS[4].t20 vss 0.08272f
C2706 BUS[4].t22 vss 0.08272f
C2707 BUS[4].n1 vss 0.44289f
C2708 BUS[4].n2 vss 0.25937f
C2709 BUS[4].t21 vss 0.08272f
C2710 BUS[4].t17 vss 0.08272f
C2711 BUS[4].n3 vss 0.44289f
C2712 BUS[4].n4 vss 0.21881f
C2713 BUS[4].t15 vss 0.66732f
C2714 BUS[4].n5 vss 0.21139f
C2715 BUS[4].t3 vss 0.08272f
C2716 BUS[4].t11 vss 0.08272f
C2717 BUS[4].n6 vss 0.44813f
C2718 BUS[4].t13 vss 0.08272f
C2719 BUS[4].t4 vss 0.08272f
C2720 BUS[4].n7 vss 0.44556f
C2721 BUS[4].n8 vss 0.25349f
C2722 BUS[4].t6 vss 0.08272f
C2723 BUS[4].t9 vss 0.08272f
C2724 BUS[4].n9 vss 0.44556f
C2725 BUS[4].n10 vss 0.14712f
C2726 BUS[4].t16 vss 0.08272f
C2727 BUS[4].t1 vss 0.08272f
C2728 BUS[4].n11 vss 0.44556f
C2729 BUS[4].n12 vss 0.14712f
C2730 BUS[4].t10 vss 0.08272f
C2731 BUS[4].t12 vss 0.08272f
C2732 BUS[4].n13 vss 0.44556f
C2733 BUS[4].n14 vss 0.14712f
C2734 BUS[4].t2 vss 0.08272f
C2735 BUS[4].t5 vss 0.08272f
C2736 BUS[4].n15 vss 0.44556f
C2737 BUS[4].n16 vss 0.14712f
C2738 BUS[4].t7 vss 0.08272f
C2739 BUS[4].t14 vss 0.08272f
C2740 BUS[4].n17 vss 0.44556f
C2741 BUS[4].n18 vss 0.14712f
C2742 BUS[4].t0 vss 0.08272f
C2743 BUS[4].t8 vss 0.08272f
C2744 BUS[4].n19 vss 0.44556f
C2745 BUS[4].n20 vss 0.11197f
C2746 BUS[4].n21 vss 0.37951f
C2747 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C2748 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C2749 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.12443f
C2750 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C2751 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C2752 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C2753 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C2754 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C2755 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C2756 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C2757 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C2758 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C2759 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C2760 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C2761 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C2762 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C2763 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C2764 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C2765 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C2766 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C2767 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C2768 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C2769 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C2770 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C2771 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C2772 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C2773 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C2774 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C2775 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C2776 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C2777 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C2778 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C2779 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C2780 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C2781 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C2782 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C2783 phi_1.t18 vss 0.12688f
C2784 phi_1.t0 vss 0.07015f
C2785 phi_1.n0 vss 0.12624f
C2786 phi_1.t4 vss 0.12688f
C2787 phi_1.t6 vss 0.07015f
C2788 phi_1.n1 vss 0.12624f
C2789 phi_1.n2 vss 1.46815f
C2790 phi_1.t8 vss 0.12688f
C2791 phi_1.t10 vss 0.07015f
C2792 phi_1.n3 vss 0.12624f
C2793 phi_1.n4 vss 1.46815f
C2794 phi_1.t16 vss 0.12688f
C2795 phi_1.t17 vss 0.07015f
C2796 phi_1.n5 vss 0.12624f
C2797 phi_1.n6 vss 1.46815f
C2798 phi_1.t19 vss 0.12688f
C2799 phi_1.t7 vss 0.07015f
C2800 phi_1.n7 vss 0.12624f
C2801 phi_1.n8 vss 1.46815f
C2802 phi_1.t11 vss 0.12688f
C2803 phi_1.t14 vss 0.07015f
C2804 phi_1.n9 vss 0.12624f
C2805 phi_1.n10 vss 1.46815f
C2806 phi_1.t12 vss 0.12688f
C2807 phi_1.t15 vss 0.07015f
C2808 phi_1.n11 vss 0.12624f
C2809 phi_1.n12 vss 1.46815f
C2810 phi_1.t1 vss 0.12688f
C2811 phi_1.t5 vss 0.07015f
C2812 phi_1.n13 vss 0.12624f
C2813 phi_1.n14 vss 1.46815f
C2814 phi_1.t9 vss 0.12688f
C2815 phi_1.t13 vss 0.07015f
C2816 phi_1.n15 vss 0.12624f
C2817 phi_1.n16 vss 1.46815f
C2818 phi_1.t2 vss 0.12688f
C2819 phi_1.t3 vss 0.07015f
C2820 phi_1.n17 vss 0.12624f
C2821 phi_1.n18 vss 1.46815f
C2822 BUS[2].t18 vss 0.08272f
C2823 BUS[2].t20 vss 0.08272f
C2824 BUS[2].n0 vss 0.44552f
C2825 BUS[2].t19 vss 0.08272f
C2826 BUS[2].t22 vss 0.08272f
C2827 BUS[2].n1 vss 0.44289f
C2828 BUS[2].n2 vss 0.25937f
C2829 BUS[2].t21 vss 0.08272f
C2830 BUS[2].t17 vss 0.08272f
C2831 BUS[2].n3 vss 0.44289f
C2832 BUS[2].n4 vss 0.21881f
C2833 BUS[2].t12 vss 0.66732f
C2834 BUS[2].n5 vss 0.21139f
C2835 BUS[2].t8 vss 0.08272f
C2836 BUS[2].t11 vss 0.08272f
C2837 BUS[2].n6 vss 0.44813f
C2838 BUS[2].t15 vss 0.08272f
C2839 BUS[2].t3 vss 0.08272f
C2840 BUS[2].n7 vss 0.44556f
C2841 BUS[2].n8 vss 0.25349f
C2842 BUS[2].t6 vss 0.08272f
C2843 BUS[2].t16 vss 0.08272f
C2844 BUS[2].n9 vss 0.44556f
C2845 BUS[2].n10 vss 0.14712f
C2846 BUS[2].t0 vss 0.08272f
C2847 BUS[2].t7 vss 0.08272f
C2848 BUS[2].n11 vss 0.44556f
C2849 BUS[2].n12 vss 0.14712f
C2850 BUS[2].t10 vss 0.08272f
C2851 BUS[2].t13 vss 0.08272f
C2852 BUS[2].n13 vss 0.44556f
C2853 BUS[2].n14 vss 0.14712f
C2854 BUS[2].t1 vss 0.08272f
C2855 BUS[2].t4 vss 0.08272f
C2856 BUS[2].n15 vss 0.44556f
C2857 BUS[2].n16 vss 0.14712f
C2858 BUS[2].t14 vss 0.08272f
C2859 BUS[2].t2 vss 0.08272f
C2860 BUS[2].n17 vss 0.44556f
C2861 BUS[2].n18 vss 0.14712f
C2862 BUS[2].t5 vss 0.08272f
C2863 BUS[2].t9 vss 0.08272f
C2864 BUS[2].n19 vss 0.44556f
C2865 BUS[2].n20 vss 0.11197f
C2866 BUS[2].n21 vss 0.37951f
C2867 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C2868 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C2869 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.12443f
C2870 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C2871 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C2872 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C2873 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C2874 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C2875 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C2876 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C2877 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C2878 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C2879 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C2880 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C2881 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C2882 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C2883 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C2884 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C2885 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C2886 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C2887 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C2888 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C2889 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C2890 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C2891 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C2892 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C2893 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C2894 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C2895 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C2896 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C2897 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C2898 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C2899 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C2900 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C2901 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C2902 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C2903 enable.t1 vss 0.01569f
C2904 enable.t7 vss 0.01886f
C2905 enable.n0 vss 0.01772f
C2906 enable.n1 vss 0.00569f
C2907 enable.t13 vss 0.01569f
C2908 enable.t0 vss 0.01886f
C2909 enable.n2 vss 0.01772f
C2910 enable.n3 vss 0.00569f
C2911 enable.t9 vss 0.01569f
C2912 enable.t15 vss 0.01886f
C2913 enable.n4 vss 0.01772f
C2914 enable.n5 vss 0.00569f
C2915 enable.t16 vss 0.01569f
C2916 enable.t5 vss 0.01886f
C2917 enable.n6 vss 0.01772f
C2918 enable.n7 vss 0.00569f
C2919 enable.t12 vss 0.01569f
C2920 enable.t19 vss 0.01886f
C2921 enable.n8 vss 0.01772f
C2922 enable.n9 vss 0.00569f
C2923 enable.t6 vss 0.01569f
C2924 enable.t17 vss 0.01886f
C2925 enable.n10 vss 0.01772f
C2926 enable.n11 vss 0.00569f
C2927 enable.t18 vss 0.01569f
C2928 enable.t8 vss 0.01886f
C2929 enable.n12 vss 0.01772f
C2930 enable.n13 vss 0.00569f
C2931 enable.t14 vss 0.01569f
C2932 enable.t4 vss 0.01886f
C2933 enable.n14 vss 0.01772f
C2934 enable.n15 vss 0.00569f
C2935 enable.t3 vss 0.01569f
C2936 enable.t11 vss 0.01886f
C2937 enable.n16 vss 0.01772f
C2938 enable.n17 vss 0.00569f
C2939 enable.t2 vss 0.01569f
C2940 enable.t10 vss 0.01886f
C2941 enable.n18 vss 0.01772f
C2942 enable.n19 vss 0.11585f
C2943 enable.n20 vss 0.1746f
C2944 enable.n21 vss 0.1746f
C2945 enable.n22 vss 0.1746f
C2946 enable.n23 vss 0.1746f
C2947 enable.n24 vss 0.1746f
C2948 enable.n25 vss 0.1746f
C2949 enable.n26 vss 0.1746f
C2950 enable.n27 vss 0.1746f
C2951 enable.n28 vss 0.1746f
C2952 BUS[10].t5 vss 0.08272f
C2953 BUS[10].t2 vss 0.08272f
C2954 BUS[10].n0 vss 0.44552f
C2955 BUS[10].t1 vss 0.08272f
C2956 BUS[10].t4 vss 0.08272f
C2957 BUS[10].n1 vss 0.44289f
C2958 BUS[10].n2 vss 0.25937f
C2959 BUS[10].t3 vss 0.08272f
C2960 BUS[10].t0 vss 0.08272f
C2961 BUS[10].n3 vss 0.44289f
C2962 BUS[10].n4 vss 0.21881f
C2963 BUS[10].t7 vss 0.66732f
C2964 BUS[10].n5 vss 0.21139f
C2965 BUS[10].t9 vss 0.08272f
C2966 BUS[10].t11 vss 0.08272f
C2967 BUS[10].n6 vss 0.44813f
C2968 BUS[10].t18 vss 0.08272f
C2969 BUS[10].t19 vss 0.08272f
C2970 BUS[10].n7 vss 0.44556f
C2971 BUS[10].n8 vss 0.25349f
C2972 BUS[10].t14 vss 0.08272f
C2973 BUS[10].t17 vss 0.08272f
C2974 BUS[10].n9 vss 0.44556f
C2975 BUS[10].n10 vss 0.14712f
C2976 BUS[10].t22 vss 0.08272f
C2977 BUS[10].t13 vss 0.08272f
C2978 BUS[10].n11 vss 0.44556f
C2979 BUS[10].n12 vss 0.14712f
C2980 BUS[10].t10 vss 0.08272f
C2981 BUS[10].t6 vss 0.08272f
C2982 BUS[10].n13 vss 0.44556f
C2983 BUS[10].n14 vss 0.14712f
C2984 BUS[10].t8 vss 0.08272f
C2985 BUS[10].t21 vss 0.08272f
C2986 BUS[10].n15 vss 0.44556f
C2987 BUS[10].n16 vss 0.14712f
C2988 BUS[10].t16 vss 0.08272f
C2989 BUS[10].t15 vss 0.08272f
C2990 BUS[10].n17 vss 0.44556f
C2991 BUS[10].n18 vss 0.14712f
C2992 BUS[10].t12 vss 0.08272f
C2993 BUS[10].t20 vss 0.08272f
C2994 BUS[10].n19 vss 0.44556f
C2995 BUS[10].n20 vss 0.11197f
C2996 BUS[10].n21 vss 0.37951f
C2997 BUS[6].t22 vss 0.08272f
C2998 BUS[6].t18 vss 0.08272f
C2999 BUS[6].n0 vss 0.44552f
C3000 BUS[6].t17 vss 0.08272f
C3001 BUS[6].t19 vss 0.08272f
C3002 BUS[6].n1 vss 0.44289f
C3003 BUS[6].n2 vss 0.25937f
C3004 BUS[6].t20 vss 0.08272f
C3005 BUS[6].t21 vss 0.08272f
C3006 BUS[6].n3 vss 0.44289f
C3007 BUS[6].n4 vss 0.21881f
C3008 BUS[6].t8 vss 0.66732f
C3009 BUS[6].n5 vss 0.21139f
C3010 BUS[6].t16 vss 0.08272f
C3011 BUS[6].t7 vss 0.08272f
C3012 BUS[6].n6 vss 0.44813f
C3013 BUS[6].t5 vss 0.08272f
C3014 BUS[6].t12 vss 0.08272f
C3015 BUS[6].n7 vss 0.44556f
C3016 BUS[6].n8 vss 0.25349f
C3017 BUS[6].t3 vss 0.08272f
C3018 BUS[6].t6 vss 0.08272f
C3019 BUS[6].n9 vss 0.44556f
C3020 BUS[6].n10 vss 0.14712f
C3021 BUS[6].t13 vss 0.08272f
C3022 BUS[6].t15 vss 0.08272f
C3023 BUS[6].n11 vss 0.44556f
C3024 BUS[6].n12 vss 0.14712f
C3025 BUS[6].t1 vss 0.08272f
C3026 BUS[6].t9 vss 0.08272f
C3027 BUS[6].n13 vss 0.44556f
C3028 BUS[6].n14 vss 0.14712f
C3029 BUS[6].t10 vss 0.08272f
C3030 BUS[6].t2 vss 0.08272f
C3031 BUS[6].n15 vss 0.44556f
C3032 BUS[6].n16 vss 0.14712f
C3033 BUS[6].t4 vss 0.08272f
C3034 BUS[6].t11 vss 0.08272f
C3035 BUS[6].n17 vss 0.44556f
C3036 BUS[6].n18 vss 0.14712f
C3037 BUS[6].t14 vss 0.08272f
C3038 BUS[6].t0 vss 0.08272f
C3039 BUS[6].n19 vss 0.44556f
C3040 BUS[6].n20 vss 0.11197f
C3041 BUS[6].n21 vss 0.37951f
C3042 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C3043 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C3044 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.12443f
C3045 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C3046 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C3047 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C3048 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C3049 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C3050 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C3051 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C3052 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C3053 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C3054 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C3055 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C3056 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C3057 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C3058 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C3059 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C3060 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C3061 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C3062 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C3063 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C3064 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C3065 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C3066 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C3067 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C3068 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C3069 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C3070 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C3071 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C3072 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C3073 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C3074 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C3075 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C3076 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C3077 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C3078 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C3079 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C3080 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.12443f
C3081 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C3082 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C3083 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C3084 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C3085 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C3086 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C3087 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C3088 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C3089 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C3090 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C3091 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C3092 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C3093 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C3094 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C3095 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C3096 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C3097 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C3098 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C3099 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C3100 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C3101 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C3102 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C3103 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C3104 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C3105 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C3106 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C3107 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C3108 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C3109 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C3110 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C3111 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C3112 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C3113 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C3114 phi_2.t18 vss 0.10942f
C3115 phi_2.t1 vss 0.0605f
C3116 phi_2.n0 vss 0.10891f
C3117 phi_2.t4 vss 0.10942f
C3118 phi_2.t11 vss 0.0605f
C3119 phi_2.n1 vss 0.10891f
C3120 phi_2.n2 vss 1.25799f
C3121 phi_2.t15 vss 0.10942f
C3122 phi_2.t17 vss 0.0605f
C3123 phi_2.n3 vss 0.10891f
C3124 phi_2.n4 vss 1.25799f
C3125 phi_2.t0 vss 0.10942f
C3126 phi_2.t3 vss 0.0605f
C3127 phi_2.n5 vss 0.10891f
C3128 phi_2.n6 vss 1.25799f
C3129 phi_2.t6 vss 0.10942f
C3130 phi_2.t7 vss 0.0605f
C3131 phi_2.n7 vss 0.10891f
C3132 phi_2.n8 vss 1.25799f
C3133 phi_2.t12 vss 0.10942f
C3134 phi_2.t14 vss 0.0605f
C3135 phi_2.n9 vss 0.10891f
C3136 phi_2.n10 vss 1.25799f
C3137 phi_2.t16 vss 0.10942f
C3138 phi_2.t5 vss 0.0605f
C3139 phi_2.n11 vss 0.10891f
C3140 phi_2.n12 vss 1.25799f
C3141 phi_2.t8 vss 0.10942f
C3142 phi_2.t10 vss 0.0605f
C3143 phi_2.n13 vss 0.10891f
C3144 phi_2.n14 vss 1.25799f
C3145 phi_2.t9 vss 0.10942f
C3146 phi_2.t13 vss 0.0605f
C3147 phi_2.n15 vss 0.10891f
C3148 phi_2.n16 vss 1.25799f
C3149 phi_2.t19 vss 0.10942f
C3150 phi_2.t2 vss 0.0605f
C3151 phi_2.n17 vss 0.10891f
C3152 phi_2.n18 vss 1.25799f
C3153 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C3154 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C3155 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.12443f
C3156 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C3157 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C3158 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C3159 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C3160 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C3161 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C3162 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C3163 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C3164 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C3165 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C3166 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C3167 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C3168 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C3169 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C3170 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C3171 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C3172 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C3173 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C3174 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C3175 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C3176 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C3177 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C3178 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C3179 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C3180 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C3181 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C3182 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C3183 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C3184 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C3185 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C3186 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C3187 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C3188 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C3189 BUS[3].t0 vss 0.08272f
C3190 BUS[3].t4 vss 0.08272f
C3191 BUS[3].n0 vss 0.44552f
C3192 BUS[3].t3 vss 0.08272f
C3193 BUS[3].t5 vss 0.08272f
C3194 BUS[3].n1 vss 0.44289f
C3195 BUS[3].n2 vss 0.25937f
C3196 BUS[3].t1 vss 0.08272f
C3197 BUS[3].t2 vss 0.08272f
C3198 BUS[3].n3 vss 0.44289f
C3199 BUS[3].n4 vss 0.21881f
C3200 BUS[3].t21 vss 0.66732f
C3201 BUS[3].n5 vss 0.21139f
C3202 BUS[3].t11 vss 0.08272f
C3203 BUS[3].t20 vss 0.08272f
C3204 BUS[3].n6 vss 0.44813f
C3205 BUS[3].t10 vss 0.08272f
C3206 BUS[3].t12 vss 0.08272f
C3207 BUS[3].n7 vss 0.44556f
C3208 BUS[3].n8 vss 0.25349f
C3209 BUS[3].t15 vss 0.08272f
C3210 BUS[3].t18 vss 0.08272f
C3211 BUS[3].n9 vss 0.44556f
C3212 BUS[3].n10 vss 0.14712f
C3213 BUS[3].t8 vss 0.08272f
C3214 BUS[3].t16 vss 0.08272f
C3215 BUS[3].n11 vss 0.44556f
C3216 BUS[3].n12 vss 0.14712f
C3217 BUS[3].t19 vss 0.08272f
C3218 BUS[3].t9 vss 0.08272f
C3219 BUS[3].n13 vss 0.44556f
C3220 BUS[3].n14 vss 0.14712f
C3221 BUS[3].t6 vss 0.08272f
C3222 BUS[3].t13 vss 0.08272f
C3223 BUS[3].n15 vss 0.44556f
C3224 BUS[3].n16 vss 0.14712f
C3225 BUS[3].t22 vss 0.08272f
C3226 BUS[3].t7 vss 0.08272f
C3227 BUS[3].n17 vss 0.44556f
C3228 BUS[3].n18 vss 0.14712f
C3229 BUS[3].t14 vss 0.08272f
C3230 BUS[3].t17 vss 0.08272f
C3231 BUS[3].n19 vss 0.44556f
C3232 BUS[3].n20 vss 0.11197f
C3233 BUS[3].n21 vss 0.37951f
C3234 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C3235 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C3236 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.12443f
C3237 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C3238 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C3239 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.1242f
C3240 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C3241 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C3242 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C3243 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C3244 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C3245 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C3246 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C3247 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C3248 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C3249 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C3250 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C3251 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C3252 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C3253 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C3254 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C3255 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C3256 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C3257 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C3258 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C3259 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C3260 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C3261 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C3262 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C3263 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C3264 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C3265 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C3266 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C3267 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C3268 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C3269 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
C3270 BUS[1].t14 vss 0.08272f
C3271 BUS[1].t15 vss 0.08272f
C3272 BUS[1].n0 vss 0.44552f
C3273 BUS[1].t16 vss 0.08272f
C3274 BUS[1].t12 vss 0.08272f
C3275 BUS[1].n1 vss 0.44289f
C3276 BUS[1].n2 vss 0.25937f
C3277 BUS[1].t17 vss 0.08272f
C3278 BUS[1].t13 vss 0.08272f
C3279 BUS[1].n3 vss 0.44289f
C3280 BUS[1].n4 vss 0.21881f
C3281 BUS[1].t22 vss 0.66732f
C3282 BUS[1].n5 vss 0.21139f
C3283 BUS[1].t2 vss 0.08272f
C3284 BUS[1].t8 vss 0.08272f
C3285 BUS[1].n6 vss 0.44813f
C3286 BUS[1].t11 vss 0.08272f
C3287 BUS[1].t1 vss 0.08272f
C3288 BUS[1].n7 vss 0.44556f
C3289 BUS[1].n8 vss 0.25349f
C3290 BUS[1].t0 vss 0.08272f
C3291 BUS[1].t10 vss 0.08272f
C3292 BUS[1].n9 vss 0.44556f
C3293 BUS[1].n10 vss 0.14712f
C3294 BUS[1].t21 vss 0.08272f
C3295 BUS[1].t19 vss 0.08272f
C3296 BUS[1].n11 vss 0.44556f
C3297 BUS[1].n12 vss 0.14712f
C3298 BUS[1].t6 vss 0.08272f
C3299 BUS[1].t4 vss 0.08272f
C3300 BUS[1].n13 vss 0.44556f
C3301 BUS[1].n14 vss 0.14712f
C3302 BUS[1].t18 vss 0.08272f
C3303 BUS[1].t5 vss 0.08272f
C3304 BUS[1].n15 vss 0.44556f
C3305 BUS[1].n16 vss 0.14712f
C3306 BUS[1].t3 vss 0.08272f
C3307 BUS[1].t9 vss 0.08272f
C3308 BUS[1].n17 vss 0.44556f
C3309 BUS[1].n18 vss 0.14712f
C3310 BUS[1].t20 vss 0.08272f
C3311 BUS[1].t7 vss 0.08272f
C3312 BUS[1].n19 vss 0.44556f
C3313 BUS[1].n20 vss 0.11197f
C3314 BUS[1].n21 vss 0.37951f
C3315 BUS[8].t2 vss 0.08272f
C3316 BUS[8].t5 vss 0.08272f
C3317 BUS[8].n0 vss 0.44552f
C3318 BUS[8].t6 vss 0.08272f
C3319 BUS[8].t7 vss 0.08272f
C3320 BUS[8].n1 vss 0.44289f
C3321 BUS[8].n2 vss 0.25937f
C3322 BUS[8].t3 vss 0.08272f
C3323 BUS[8].t4 vss 0.08272f
C3324 BUS[8].n3 vss 0.44289f
C3325 BUS[8].n4 vss 0.21881f
C3326 BUS[8].t10 vss 0.66732f
C3327 BUS[8].n5 vss 0.21139f
C3328 BUS[8].t8 vss 0.08272f
C3329 BUS[8].t0 vss 0.08272f
C3330 BUS[8].n6 vss 0.44813f
C3331 BUS[8].t19 vss 0.08272f
C3332 BUS[8].t15 vss 0.08272f
C3333 BUS[8].n7 vss 0.44556f
C3334 BUS[8].n8 vss 0.25349f
C3335 BUS[8].t22 vss 0.08272f
C3336 BUS[8].t16 vss 0.08272f
C3337 BUS[8].n9 vss 0.44556f
C3338 BUS[8].n10 vss 0.14712f
C3339 BUS[8].t21 vss 0.08272f
C3340 BUS[8].t18 vss 0.08272f
C3341 BUS[8].n11 vss 0.44556f
C3342 BUS[8].n12 vss 0.14712f
C3343 BUS[8].t1 vss 0.08272f
C3344 BUS[8].t20 vss 0.08272f
C3345 BUS[8].n13 vss 0.44556f
C3346 BUS[8].n14 vss 0.14712f
C3347 BUS[8].t9 vss 0.08272f
C3348 BUS[8].t14 vss 0.08272f
C3349 BUS[8].n15 vss 0.44556f
C3350 BUS[8].n16 vss 0.14712f
C3351 BUS[8].t12 vss 0.08272f
C3352 BUS[8].t11 vss 0.08272f
C3353 BUS[8].n17 vss 0.44556f
C3354 BUS[8].n18 vss 0.14712f
C3355 BUS[8].t13 vss 0.08272f
C3356 BUS[8].t17 vss 0.08272f
C3357 BUS[8].n19 vss 0.44556f
C3358 BUS[8].n20 vss 0.11197f
C3359 BUS[8].n21 vss 0.37951f
C3360 vdd.t8 vss 0.0089f
C3361 vdd.t497 vss 0.00436f
C3362 vdd.n0 vss 0.01891f
C3363 vdd.t517 vss 0.0111f
C3364 vdd.t130 vss 0.00591f
C3365 vdd.t453 vss 0.00591f
C3366 vdd.n1 vss 0.01262f
C3367 vdd.t128 vss 0.02243f
C3368 vdd.t496 vss 0.10168f
C3369 vdd.t7 vss 0.16586f
C3370 vdd.t516 vss 0.13628f
C3371 vdd.t6 vss 0.09296f
C3372 vdd.t465 vss 0.11726f
C3373 vdd.t452 vss 0.11726f
C3374 vdd.t129 vss 0.16691f
C3375 vdd.t127 vss 0.1928f
C3376 vdd.n2 vss 0.12094f
C3377 vdd.t99 vss 0.0089f
C3378 vdd.t243 vss 0.00436f
C3379 vdd.n3 vss 0.01891f
C3380 vdd.t451 vss 0.0111f
C3381 vdd.t270 vss 0.00591f
C3382 vdd.t413 vss 0.00591f
C3383 vdd.n4 vss 0.01262f
C3384 vdd.t272 vss 0.02243f
C3385 vdd.t449 vss 0.01933f
C3386 vdd.t22 vss 0.01907f
C3387 vdd.t173 vss 0.02206f
C3388 vdd.t242 vss 0.10168f
C3389 vdd.t98 vss 0.16586f
C3390 vdd.t450 vss 0.13628f
C3391 vdd.t97 vss 0.09296f
C3392 vdd.t215 vss 0.11726f
C3393 vdd.t412 vss 0.11726f
C3394 vdd.t269 vss 0.16691f
C3395 vdd.t271 vss 0.18249f
C3396 vdd.t448 vss 0.08187f
C3397 vdd.t21 vss 0.1199f
C3398 vdd.t172 vss 0.12862f
C3399 vdd.n5 vss 0.16821f
C3400 vdd.n6 vss 0.12147f
C3401 vdd.t369 vss 0.0089f
C3402 vdd.t529 vss 0.00436f
C3403 vdd.n7 vss 0.01891f
C3404 vdd.t447 vss 0.0111f
C3405 vdd.t241 vss 0.00591f
C3406 vdd.t222 vss 0.00591f
C3407 vdd.n8 vss 0.01262f
C3408 vdd.t239 vss 0.02243f
C3409 vdd.t528 vss 0.10168f
C3410 vdd.t368 vss 0.16586f
C3411 vdd.t446 vss 0.13628f
C3412 vdd.t370 vss 0.09296f
C3413 vdd.t136 vss 0.11726f
C3414 vdd.t221 vss 0.11726f
C3415 vdd.t240 vss 0.16691f
C3416 vdd.t238 vss 0.1928f
C3417 vdd.n9 vss 0.12094f
C3418 vdd.t421 vss 0.0089f
C3419 vdd.t255 vss 0.00436f
C3420 vdd.n10 vss 0.01891f
C3421 vdd.t52 vss 0.0111f
C3422 vdd.t175 vss 0.00591f
C3423 vdd.t192 vss 0.00591f
C3424 vdd.n11 vss 0.01262f
C3425 vdd.t177 vss 0.02243f
C3426 vdd.t41 vss 0.01933f
C3427 vdd.t460 vss 0.01907f
C3428 vdd.t65 vss 0.02206f
C3429 vdd.t254 vss 0.10168f
C3430 vdd.t420 vss 0.16586f
C3431 vdd.t51 vss 0.13628f
C3432 vdd.t419 vss 0.09296f
C3433 vdd.t212 vss 0.11726f
C3434 vdd.t191 vss 0.11726f
C3435 vdd.t174 vss 0.16691f
C3436 vdd.t176 vss 0.18249f
C3437 vdd.t40 vss 0.08187f
C3438 vdd.t459 vss 0.1199f
C3439 vdd.t64 vss 0.12862f
C3440 vdd.n12 vss 0.16821f
C3441 vdd.n13 vss 0.12147f
C3442 vdd.t60 vss 0.0089f
C3443 vdd.t495 vss 0.00436f
C3444 vdd.n14 vss 0.01891f
C3445 vdd.t39 vss 0.0111f
C3446 vdd.t29 vss 0.00591f
C3447 vdd.t488 vss 0.00591f
C3448 vdd.n15 vss 0.01262f
C3449 vdd.t31 vss 0.02243f
C3450 vdd.t494 vss 0.10168f
C3451 vdd.t59 vss 0.16586f
C3452 vdd.t38 vss 0.13628f
C3453 vdd.t61 vss 0.09296f
C3454 vdd.t515 vss 0.11726f
C3455 vdd.t487 vss 0.11726f
C3456 vdd.t28 vss 0.16691f
C3457 vdd.t30 vss 0.1928f
C3458 vdd.n16 vss 0.12094f
C3459 vdd.t330 vss 0.0089f
C3460 vdd.t253 vss 0.00436f
C3461 vdd.n17 vss 0.01891f
C3462 vdd.t471 vss 0.0111f
C3463 vdd.t122 vss 0.00591f
C3464 vdd.t135 vss 0.00591f
C3465 vdd.n18 vss 0.01262f
C3466 vdd.t124 vss 0.02243f
C3467 vdd.t510 vss 0.01933f
C3468 vdd.t477 vss 0.01907f
C3469 vdd.t120 vss 0.02206f
C3470 vdd.t252 vss 0.10168f
C3471 vdd.t329 vss 0.16586f
C3472 vdd.t470 vss 0.13628f
C3473 vdd.t328 vss 0.09296f
C3474 vdd.t137 vss 0.11726f
C3475 vdd.t134 vss 0.11726f
C3476 vdd.t121 vss 0.16691f
C3477 vdd.t123 vss 0.18249f
C3478 vdd.t509 vss 0.08187f
C3479 vdd.t476 vss 0.1199f
C3480 vdd.t119 vss 0.12862f
C3481 vdd.n19 vss 0.16821f
C3482 vdd.n20 vss 0.12147f
C3483 vdd.t160 vss 0.0089f
C3484 vdd.t69 vss 0.00436f
C3485 vdd.n21 vss 0.01891f
C3486 vdd.t512 vss 0.0111f
C3487 vdd.t92 vss 0.00591f
C3488 vdd.t503 vss 0.00591f
C3489 vdd.n22 vss 0.01262f
C3490 vdd.t90 vss 0.02243f
C3491 vdd.t68 vss 0.10168f
C3492 vdd.t159 vss 0.16586f
C3493 vdd.t511 vss 0.13628f
C3494 vdd.t158 vss 0.09296f
C3495 vdd.t110 vss 0.11726f
C3496 vdd.t502 vss 0.11726f
C3497 vdd.t91 vss 0.16691f
C3498 vdd.t89 vss 0.1928f
C3499 vdd.n23 vss 0.12094f
C3500 vdd.t260 vss 0.0089f
C3501 vdd.t35 vss 0.00436f
C3502 vdd.n24 vss 0.01891f
C3503 vdd.t171 vss 0.0111f
C3504 vdd.t54 vss 0.00591f
C3505 vdd.t162 vss 0.00591f
C3506 vdd.n25 vss 0.01262f
C3507 vdd.t56 vss 0.02243f
C3508 vdd.t268 vss 0.01933f
C3509 vdd.t469 vss 0.01907f
C3510 vdd.t112 vss 0.02206f
C3511 vdd.t34 vss 0.10168f
C3512 vdd.t259 vss 0.16586f
C3513 vdd.t170 vss 0.13628f
C3514 vdd.t258 vss 0.09296f
C3515 vdd.t180 vss 0.11726f
C3516 vdd.t161 vss 0.11726f
C3517 vdd.t53 vss 0.16691f
C3518 vdd.t55 vss 0.18249f
C3519 vdd.t267 vss 0.08187f
C3520 vdd.t468 vss 0.1199f
C3521 vdd.t111 vss 0.12862f
C3522 vdd.n26 vss 0.16821f
C3523 vdd.n27 vss 0.12147f
C3524 vdd.t417 vss 0.0089f
C3525 vdd.t67 vss 0.00436f
C3526 vdd.n28 vss 0.01891f
C3527 vdd.t266 vss 0.0111f
C3528 vdd.t424 vss 0.00591f
C3529 vdd.t492 vss 0.00591f
C3530 vdd.n29 vss 0.01262f
C3531 vdd.t426 vss 0.02243f
C3532 vdd.t66 vss 0.10168f
C3533 vdd.t416 vss 0.16586f
C3534 vdd.t265 vss 0.13628f
C3535 vdd.t418 vss 0.09296f
C3536 vdd.t391 vss 0.11726f
C3537 vdd.t491 vss 0.11726f
C3538 vdd.t423 vss 0.16691f
C3539 vdd.t425 vss 0.1928f
C3540 vdd.n30 vss 0.12094f
C3541 vdd.t132 vss 0.0089f
C3542 vdd.t290 vss 0.00436f
C3543 vdd.n31 vss 0.01891f
C3544 vdd.t209 vss 0.0111f
C3545 vdd.t362 vss 0.00591f
C3546 vdd.t96 vss 0.00591f
C3547 vdd.n32 vss 0.01262f
C3548 vdd.t364 vss 0.02243f
C3549 vdd.t157 vss 0.01933f
C3550 vdd.t458 vss 0.01907f
C3551 vdd.t126 vss 0.02206f
C3552 vdd.t289 vss 0.10168f
C3553 vdd.t131 vss 0.16586f
C3554 vdd.t208 vss 0.13628f
C3555 vdd.t133 vss 0.09296f
C3556 vdd.t62 vss 0.11726f
C3557 vdd.t95 vss 0.11726f
C3558 vdd.t361 vss 0.16691f
C3559 vdd.t363 vss 0.18249f
C3560 vdd.t156 vss 0.08187f
C3561 vdd.t457 vss 0.1199f
C3562 vdd.t125 vss 0.12862f
C3563 vdd.n33 vss 0.16821f
C3564 vdd.n34 vss 0.12147f
C3565 vdd.t139 vss 0.0089f
C3566 vdd.t257 vss 0.00436f
C3567 vdd.n35 vss 0.01891f
C3568 vdd.t155 vss 0.0111f
C3569 vdd.t376 vss 0.00591f
C3570 vdd.t337 vss 0.00591f
C3571 vdd.n36 vss 0.01262f
C3572 vdd.t378 vss 0.02243f
C3573 vdd.t256 vss 0.10168f
C3574 vdd.t138 vss 0.16586f
C3575 vdd.t154 vss 0.13628f
C3576 vdd.t140 vss 0.09296f
C3577 vdd.t338 vss 0.11726f
C3578 vdd.t336 vss 0.11726f
C3579 vdd.t375 vss 0.16691f
C3580 vdd.t377 vss 0.1928f
C3581 vdd.n37 vss 0.12094f
C3582 vdd.t190 vss 0.0089f
C3583 vdd.t346 vss 0.00436f
C3584 vdd.n38 vss 0.01891f
C3585 vdd.t402 vss 0.0111f
C3586 vdd.t479 vss 0.00591f
C3587 vdd.t94 vss 0.00591f
C3588 vdd.n39 vss 0.01262f
C3589 vdd.t481 vss 0.02243f
C3590 vdd.t292 vss 0.01933f
C3591 vdd.t20 vss 0.01907f
C3592 vdd.t382 vss 0.02206f
C3593 vdd.t345 vss 0.10168f
C3594 vdd.t189 vss 0.16586f
C3595 vdd.t401 vss 0.13628f
C3596 vdd.t188 vss 0.09296f
C3597 vdd.t429 vss 0.11726f
C3598 vdd.t93 vss 0.11726f
C3599 vdd.t478 vss 0.16691f
C3600 vdd.t480 vss 0.18249f
C3601 vdd.t291 vss 0.08187f
C3602 vdd.t19 vss 0.1199f
C3603 vdd.t381 vss 0.12862f
C3604 vdd.n40 vss 0.16821f
C3605 vdd.n41 vss 0.12147f
C3606 vdd.t334 vss 0.0089f
C3607 vdd.t301 vss 0.00436f
C3608 vdd.n42 vss 0.01891f
C3609 vdd.t294 vss 0.0111f
C3610 vdd.t166 vss 0.00591f
C3611 vdd.t372 vss 0.00591f
C3612 vdd.n43 vss 0.01262f
C3613 vdd.t164 vss 0.02243f
C3614 vdd.t300 vss 0.10168f
C3615 vdd.t333 vss 0.16586f
C3616 vdd.t293 vss 0.13628f
C3617 vdd.t335 vss 0.09296f
C3618 vdd.t169 vss 0.11726f
C3619 vdd.t371 vss 0.11726f
C3620 vdd.t165 vss 0.16691f
C3621 vdd.t163 vss 0.1928f
C3622 vdd.n44 vss 0.12094f
C3623 vdd.t406 vss 0.0089f
C3624 vdd.t146 vss 0.00436f
C3625 vdd.n45 vss 0.01891f
C3626 vdd.t179 vss 0.0111f
C3627 vdd.t400 vss 0.00591f
C3628 vdd.t332 vss 0.00591f
C3629 vdd.n46 vss 0.01262f
C3630 vdd.t398 vss 0.02243f
C3631 vdd.t390 vss 0.01933f
C3632 vdd.t483 vss 0.01907f
C3633 vdd.t506 vss 0.02206f
C3634 vdd.t145 vss 0.10168f
C3635 vdd.t405 vss 0.16586f
C3636 vdd.t178 vss 0.13628f
C3637 vdd.t404 vss 0.09296f
C3638 vdd.t23 vss 0.11726f
C3639 vdd.t331 vss 0.11726f
C3640 vdd.t399 vss 0.16691f
C3641 vdd.t397 vss 0.18249f
C3642 vdd.t389 vss 0.08187f
C3643 vdd.t482 vss 0.1199f
C3644 vdd.t505 vss 0.12862f
C3645 vdd.n47 vss 0.16821f
C3646 vdd.n48 vss 0.12147f
C3647 vdd.t148 vss 0.0089f
C3648 vdd.t527 vss 0.00436f
C3649 vdd.n49 vss 0.01891f
C3650 vdd.t388 vss 0.0111f
C3651 vdd.t18 vss 0.00591f
C3652 vdd.t251 vss 0.00591f
C3653 vdd.n50 vss 0.01262f
C3654 vdd.t16 vss 0.02243f
C3655 vdd.t526 vss 0.10168f
C3656 vdd.t147 vss 0.16586f
C3657 vdd.t387 vss 0.13628f
C3658 vdd.t149 vss 0.09296f
C3659 vdd.t63 vss 0.11726f
C3660 vdd.t250 vss 0.11726f
C3661 vdd.t17 vss 0.16691f
C3662 vdd.t15 vss 0.1928f
C3663 vdd.n51 vss 0.12094f
C3664 vdd.t436 vss 0.0089f
C3665 vdd.t33 vss 0.00436f
C3666 vdd.n52 vss 0.01891f
C3667 vdd.t182 vss 0.0111f
C3668 vdd.t207 vss 0.00591f
C3669 vdd.t307 vss 0.00591f
C3670 vdd.n53 vss 0.01262f
C3671 vdd.t205 vss 0.02243f
C3672 vdd.t443 vss 0.01933f
C3673 vdd.t467 vss 0.01907f
C3674 vdd.t428 vss 0.02206f
C3675 vdd.t32 vss 0.10168f
C3676 vdd.t435 vss 0.16586f
C3677 vdd.t181 vss 0.13628f
C3678 vdd.t437 vss 0.09296f
C3679 vdd.t486 vss 0.11726f
C3680 vdd.t306 vss 0.11726f
C3681 vdd.t206 vss 0.16691f
C3682 vdd.t204 vss 0.18249f
C3683 vdd.t442 vss 0.08187f
C3684 vdd.t466 vss 0.1199f
C3685 vdd.t427 vss 0.12862f
C3686 vdd.n54 vss 0.16821f
C3687 vdd.n55 vss 0.12147f
C3688 vdd.t144 vss 0.0089f
C3689 vdd.t445 vss 0.00436f
C3690 vdd.n56 vss 0.01891f
C3691 vdd.t441 vss 0.0111f
C3692 vdd.t197 vss 0.00591f
C3693 vdd.t71 vss 0.00591f
C3694 vdd.n57 vss 0.01262f
C3695 vdd.t199 vss 0.02243f
C3696 vdd.t444 vss 0.10168f
C3697 vdd.t143 vss 0.16586f
C3698 vdd.t440 vss 0.13628f
C3699 vdd.t142 vss 0.09296f
C3700 vdd.t141 vss 0.11726f
C3701 vdd.t70 vss 0.11726f
C3702 vdd.t196 vss 0.16691f
C3703 vdd.t198 vss 0.1928f
C3704 vdd.n58 vss 0.12094f
C3705 vdd.t279 vss 0.0089f
C3706 vdd.t344 vss 0.00436f
C3707 vdd.n59 vss 0.01891f
C3708 vdd.t201 vss 0.0111f
C3709 vdd.t384 vss 0.00591f
C3710 vdd.t58 vss 0.00591f
C3711 vdd.n60 vss 0.01262f
C3712 vdd.t386 vss 0.02243f
C3713 vdd.t12 vss 0.01933f
C3714 vdd.t464 vss 0.01907f
C3715 vdd.t168 vss 0.02206f
C3716 vdd.t343 vss 0.10168f
C3717 vdd.t278 vss 0.16586f
C3718 vdd.t200 vss 0.13628f
C3719 vdd.t280 vss 0.09296f
C3720 vdd.t403 vss 0.11726f
C3721 vdd.t57 vss 0.11726f
C3722 vdd.t383 vss 0.16691f
C3723 vdd.t385 vss 0.18249f
C3724 vdd.t11 vss 0.08187f
C3725 vdd.t463 vss 0.1199f
C3726 vdd.t167 vss 0.12862f
C3727 vdd.n61 vss 0.16821f
C3728 vdd.n62 vss 0.12147f
C3729 vdd.t475 vss 0.0089f
C3730 vdd.t303 vss 0.00436f
C3731 vdd.n63 vss 0.01891f
C3732 vdd.t10 vss 0.0111f
C3733 vdd.t103 vss 0.00591f
C3734 vdd.t211 vss 0.00591f
C3735 vdd.n64 vss 0.01262f
C3736 vdd.t101 vss 0.02243f
C3737 vdd.t302 vss 0.10168f
C3738 vdd.t474 vss 0.16586f
C3739 vdd.t9 vss 0.13628f
C3740 vdd.t473 vss 0.09296f
C3741 vdd.t472 vss 0.11726f
C3742 vdd.t210 vss 0.11726f
C3743 vdd.t102 vss 0.16691f
C3744 vdd.t100 vss 0.1928f
C3745 vdd.n65 vss 0.12094f
C3746 vdd.t434 vss 0.0089f
C3747 vdd.t37 vss 0.00436f
C3748 vdd.n66 vss 0.01891f
C3749 vdd.t501 vss 0.0111f
C3750 vdd.t217 vss 0.00591f
C3751 vdd.t524 vss 0.00591f
C3752 vdd.n67 vss 0.01262f
C3753 vdd.t219 vss 0.02243f
C3754 vdd.t341 vss 0.01933f
C3755 vdd.t462 vss 0.01907f
C3756 vdd.t411 vss 0.02206f
C3757 vdd.t36 vss 0.10168f
C3758 vdd.t433 vss 0.16586f
C3759 vdd.t500 vss 0.13628f
C3760 vdd.t432 vss 0.09296f
C3761 vdd.t456 vss 0.11726f
C3762 vdd.t523 vss 0.11726f
C3763 vdd.t216 vss 0.16691f
C3764 vdd.t218 vss 0.18249f
C3765 vdd.t340 vss 0.08187f
C3766 vdd.t461 vss 0.1199f
C3767 vdd.t410 vss 0.13029f
C3768 vdd.n68 vss 0.33568f
C3769 vdd.n69 vss 0.05099f
C3770 vdd.n70 vss 0.05384f
C3771 vdd.n71 vss 0.07323f
C3772 vdd.n72 vss 0.11512f
C3773 vdd.n73 vss 0.10389f
C3774 vdd.n74 vss 0.07151f
C3775 vdd.n75 vss 0.06428f
C3776 vdd.n76 vss 0.07553f
C3777 vdd.n77 vss 0.11512f
C3778 vdd.n78 vss 0.10389f
C3779 vdd.n79 vss 0.0506f
C3780 vdd.n80 vss 0.05123f
C3781 vdd.n81 vss 0.06413f
C3782 vdd.n82 vss 0.05917f
C3783 vdd.n83 vss 0.05099f
C3784 vdd.n84 vss 0.05384f
C3785 vdd.n85 vss 0.07323f
C3786 vdd.n86 vss 0.11512f
C3787 vdd.n87 vss 0.10389f
C3788 vdd.n88 vss 0.07151f
C3789 vdd.n89 vss 0.06428f
C3790 vdd.n90 vss 0.07553f
C3791 vdd.n91 vss 0.11512f
C3792 vdd.n92 vss 0.10389f
C3793 vdd.n93 vss 0.0506f
C3794 vdd.n94 vss 0.05123f
C3795 vdd.n95 vss 0.06413f
C3796 vdd.n96 vss 0.05917f
C3797 vdd.n97 vss 0.05099f
C3798 vdd.n98 vss 0.05384f
C3799 vdd.n99 vss 0.07323f
C3800 vdd.n100 vss 0.11512f
C3801 vdd.n101 vss 0.10389f
C3802 vdd.n102 vss 0.07151f
C3803 vdd.n103 vss 0.06428f
C3804 vdd.n104 vss 0.07553f
C3805 vdd.n105 vss 0.11512f
C3806 vdd.n106 vss 0.10389f
C3807 vdd.n107 vss 0.0506f
C3808 vdd.n108 vss 0.05123f
C3809 vdd.n109 vss 0.06413f
C3810 vdd.n110 vss 0.05917f
C3811 vdd.n111 vss 0.05099f
C3812 vdd.n112 vss 0.05384f
C3813 vdd.n113 vss 0.07323f
C3814 vdd.n114 vss 0.11512f
C3815 vdd.n115 vss 0.10389f
C3816 vdd.n116 vss 0.07151f
C3817 vdd.n117 vss 0.06428f
C3818 vdd.n118 vss 0.07553f
C3819 vdd.n119 vss 0.11512f
C3820 vdd.n120 vss 0.10389f
C3821 vdd.n121 vss 0.0506f
C3822 vdd.n122 vss 0.05123f
C3823 vdd.n123 vss 0.06413f
C3824 vdd.n124 vss 0.05917f
C3825 vdd.n125 vss 0.05099f
C3826 vdd.n126 vss 0.05384f
C3827 vdd.n127 vss 0.07323f
C3828 vdd.n128 vss 0.11512f
C3829 vdd.n129 vss 0.10389f
C3830 vdd.n130 vss 0.07151f
C3831 vdd.n131 vss 0.06428f
C3832 vdd.n132 vss 0.07553f
C3833 vdd.n133 vss 0.11512f
C3834 vdd.n134 vss 0.10389f
C3835 vdd.n135 vss 0.0506f
C3836 vdd.n136 vss 0.05123f
C3837 vdd.n137 vss 0.06413f
C3838 vdd.n138 vss 0.05917f
C3839 vdd.n139 vss 0.05099f
C3840 vdd.n140 vss 0.05384f
C3841 vdd.n141 vss 0.07323f
C3842 vdd.n142 vss 0.11512f
C3843 vdd.n143 vss 0.10389f
C3844 vdd.n144 vss 0.07151f
C3845 vdd.n145 vss 0.06428f
C3846 vdd.n146 vss 0.07553f
C3847 vdd.n147 vss 0.11512f
C3848 vdd.n148 vss 0.10389f
C3849 vdd.n149 vss 0.0506f
C3850 vdd.n150 vss 0.05123f
C3851 vdd.n151 vss 0.06413f
C3852 vdd.n152 vss 0.05917f
C3853 vdd.n153 vss 0.05099f
C3854 vdd.n154 vss 0.05384f
C3855 vdd.n155 vss 0.07323f
C3856 vdd.n156 vss 0.11512f
C3857 vdd.n157 vss 0.10389f
C3858 vdd.n158 vss 0.07151f
C3859 vdd.n159 vss 0.06428f
C3860 vdd.n160 vss 0.07553f
C3861 vdd.n161 vss 0.11512f
C3862 vdd.n162 vss 0.10389f
C3863 vdd.n163 vss 0.0506f
C3864 vdd.n164 vss 0.05123f
C3865 vdd.n165 vss 0.06413f
C3866 vdd.n166 vss 0.05917f
C3867 vdd.n167 vss 0.05099f
C3868 vdd.n168 vss 0.05384f
C3869 vdd.n169 vss 0.07323f
C3870 vdd.n170 vss 0.11512f
C3871 vdd.n171 vss 0.10389f
C3872 vdd.n172 vss 0.07151f
C3873 vdd.n173 vss 0.06428f
C3874 vdd.n174 vss 0.07553f
C3875 vdd.n175 vss 0.11512f
C3876 vdd.n176 vss 0.10389f
C3877 vdd.n177 vss 0.0506f
C3878 vdd.n178 vss 0.05123f
C3879 vdd.n179 vss 0.06413f
C3880 vdd.n180 vss 0.05917f
C3881 vdd.n181 vss 0.05099f
C3882 vdd.n182 vss 0.05384f
C3883 vdd.n183 vss 0.07323f
C3884 vdd.n184 vss 0.11512f
C3885 vdd.n185 vss 0.10389f
C3886 vdd.n186 vss 0.07151f
C3887 vdd.n187 vss 0.06428f
C3888 vdd.n188 vss 0.07553f
C3889 vdd.n189 vss 0.11512f
C3890 vdd.n190 vss 0.10389f
C3891 vdd.n191 vss 0.0506f
C3892 vdd.n192 vss 0.05123f
C3893 vdd.n193 vss 0.06413f
C3894 vdd.n194 vss 0.05917f
C3895 vdd.n195 vss 0.05099f
C3896 vdd.n196 vss 0.05384f
C3897 vdd.n197 vss 0.07323f
C3898 vdd.n198 vss 0.11512f
C3899 vdd.n199 vss 0.10389f
C3900 vdd.n200 vss 0.07151f
C3901 vdd.n201 vss 0.06428f
C3902 vdd.n202 vss 0.07553f
C3903 vdd.n203 vss 0.11512f
C3904 vdd.n204 vss 0.10389f
C3905 vdd.n205 vss 0.0506f
C3906 vdd.n206 vss 0.19265f
C3907 vdd.t454 vss 0.17868f
C3908 vdd.t455 vss 0.02206f
C3909 vdd.t522 vss 0.33339f
C3910 vdd.t227 vss 0.14187f
C3911 vdd.t520 vss 0.14187f
C3912 vdd.t286 vss 0.14187f
C3913 vdd.t108 vss 0.14187f
C3914 vdd.t225 vss 0.14187f
C3915 vdd.t518 vss 0.14187f
C3916 vdd.t109 vss 0.14187f
C3917 vdd.t226 vss 0.14187f
C3918 vdd.t519 vss 0.14187f
C3919 vdd.t521 vss 0.14187f
C3920 vdd.t287 vss 0.14187f
C3921 vdd.t42 vss 0.14187f
C3922 vdd.t43 vss 0.14187f
C3923 vdd.t288 vss 0.14187f
C3924 vdd.t228 vss 0.14187f
C3925 vdd.t44 vss 0.18766f
C3926 vdd.t152 vss 0.17868f
C3927 vdd.t153 vss 0.02206f
C3928 vdd.t2 vss 0.33339f
C3929 vdd.t5 vss 0.14187f
C3930 vdd.t105 vss 0.14187f
C3931 vdd.t193 vss 0.14187f
C3932 vdd.t0 vss 0.14187f
C3933 vdd.t24 vss 0.14187f
C3934 vdd.t194 vss 0.14187f
C3935 vdd.t1 vss 0.14187f
C3936 vdd.t4 vss 0.14187f
C3937 vdd.t118 vss 0.14187f
C3938 vdd.t220 vss 0.14187f
C3939 vdd.t507 vss 0.14187f
C3940 vdd.t104 vss 0.14187f
C3941 vdd.t25 vss 0.14187f
C3942 vdd.t195 vss 0.14187f
C3943 vdd.t3 vss 0.14187f
C3944 vdd.t117 vss 0.18766f
C3945 vdd.t379 vss 0.17868f
C3946 vdd.t380 vss 0.02206f
C3947 vdd.t114 vss 0.33339f
C3948 vdd.t229 vss 0.14187f
C3949 vdd.t430 vss 0.14187f
C3950 vdd.t235 vss 0.14187f
C3951 vdd.t113 vss 0.14187f
C3952 vdd.t431 vss 0.14187f
C3953 vdd.t184 vss 0.14187f
C3954 vdd.t233 vss 0.14187f
C3955 vdd.t46 vss 0.14187f
C3956 vdd.t230 vss 0.14187f
C3957 vdd.t234 vss 0.14187f
C3958 vdd.t47 vss 0.14187f
C3959 vdd.t231 vss 0.14187f
C3960 vdd.t247 vss 0.14187f
C3961 vdd.t249 vss 0.14187f
C3962 vdd.t45 vss 0.14187f
C3963 vdd.t248 vss 0.18766f
C3964 vdd.t484 vss 0.17868f
C3965 vdd.t485 vss 0.02206f
C3966 vdd.t322 vss 0.33339f
C3967 vdd.t308 vss 0.14187f
C3968 vdd.t264 vss 0.14187f
C3969 vdd.t323 vss 0.14187f
C3970 vdd.t309 vss 0.14187f
C3971 vdd.t312 vss 0.14187f
C3972 vdd.t374 vss 0.14187f
C3973 vdd.t311 vss 0.14187f
C3974 vdd.t438 vss 0.14187f
C3975 vdd.t321 vss 0.14187f
C3976 vdd.t356 vss 0.14187f
C3977 vdd.t439 vss 0.14187f
C3978 vdd.t183 vss 0.14187f
C3979 vdd.t313 vss 0.14187f
C3980 vdd.t310 vss 0.14187f
C3981 vdd.t320 vss 0.14187f
C3982 vdd.t373 vss 0.18766f
C3983 vdd.t150 vss 0.17868f
C3984 vdd.t151 vss 0.02206f
C3985 vdd.t83 vss 0.33339f
C3986 vdd.t81 vss 0.14187f
C3987 vdd.t73 vss 0.14187f
C3988 vdd.t82 vss 0.14187f
C3989 vdd.t85 vss 0.14187f
C3990 vdd.t78 vss 0.14187f
C3991 vdd.t75 vss 0.14187f
C3992 vdd.t84 vss 0.14187f
C3993 vdd.t77 vss 0.14187f
C3994 vdd.t74 vss 0.14187f
C3995 vdd.t72 vss 0.14187f
C3996 vdd.t87 vss 0.14187f
C3997 vdd.t80 vss 0.14187f
C3998 vdd.t88 vss 0.14187f
C3999 vdd.t86 vss 0.14187f
C4000 vdd.t79 vss 0.14187f
C4001 vdd.t76 vss 0.18766f
C4002 vdd.t392 vss 0.17868f
C4003 vdd.t393 vss 0.02206f
C4004 vdd.t237 vss 0.33339f
C4005 vdd.t285 vss 0.14187f
C4006 vdd.t350 vss 0.14187f
C4007 vdd.t49 vss 0.14187f
C4008 vdd.t394 vss 0.14187f
C4009 vdd.t396 vss 0.14187f
C4010 vdd.t50 vss 0.14187f
C4011 vdd.t236 vss 0.14187f
C4012 vdd.t284 vss 0.14187f
C4013 vdd.t349 vss 0.14187f
C4014 vdd.t351 vss 0.14187f
C4015 vdd.t245 vss 0.14187f
C4016 vdd.t395 vss 0.14187f
C4017 vdd.t48 vss 0.14187f
C4018 vdd.t246 vss 0.14187f
C4019 vdd.t244 vss 0.14187f
C4020 vdd.t493 vss 0.18766f
C4021 vdd.t498 vss 0.17868f
C4022 vdd.t499 vss 0.02206f
C4023 vdd.t325 vss 0.33339f
C4024 vdd.t297 vss 0.14187f
C4025 vdd.t274 vss 0.14187f
C4026 vdd.t513 vss 0.14187f
C4027 vdd.t504 vss 0.14187f
C4028 vdd.t275 vss 0.14187f
C4029 vdd.t514 vss 0.14187f
C4030 vdd.t342 vss 0.14187f
C4031 vdd.t348 vss 0.14187f
C4032 vdd.t316 vss 0.14187f
C4033 vdd.t347 vss 0.14187f
C4034 vdd.t296 vss 0.14187f
C4035 vdd.t317 vss 0.14187f
C4036 vdd.t232 vss 0.14187f
C4037 vdd.t324 vss 0.14187f
C4038 vdd.t366 vss 0.14187f
C4039 vdd.t304 vss 0.18766f
C4040 vdd.t26 vss 0.17868f
C4041 vdd.t27 vss 0.02206f
C4042 vdd.t185 vss 0.33339f
C4043 vdd.t282 vss 0.14187f
C4044 vdd.t261 vss 0.14187f
C4045 vdd.t186 vss 0.14187f
C4046 vdd.t187 vss 0.14187f
C4047 vdd.t262 vss 0.14187f
C4048 vdd.t116 vss 0.14187f
C4049 vdd.t408 vss 0.14187f
C4050 vdd.t14 vss 0.14187f
C4051 vdd.t283 vss 0.14187f
C4052 vdd.t409 vss 0.14187f
C4053 vdd.t281 vss 0.14187f
C4054 vdd.t525 vss 0.14187f
C4055 vdd.t263 vss 0.14187f
C4056 vdd.t407 vss 0.14187f
C4057 vdd.t13 vss 0.14187f
C4058 vdd.t115 vss 0.18766f
C4059 vdd.t489 vss 0.17868f
C4060 vdd.t490 vss 0.02206f
C4061 vdd.t315 vss 0.33339f
C4062 vdd.t415 vss 0.14187f
C4063 vdd.t365 vss 0.14187f
C4064 vdd.t273 vss 0.14187f
C4065 vdd.t299 vss 0.14187f
C4066 vdd.t203 vss 0.14187f
C4067 vdd.t352 vss 0.14187f
C4068 vdd.t508 vss 0.14187f
C4069 vdd.t414 vss 0.14187f
C4070 vdd.t353 vss 0.14187f
C4071 vdd.t314 vss 0.14187f
C4072 vdd.t339 vss 0.14187f
C4073 vdd.t295 vss 0.14187f
C4074 vdd.t357 vss 0.14187f
C4075 vdd.t298 vss 0.14187f
C4076 vdd.t202 vss 0.14187f
C4077 vdd.t358 vss 0.18766f
C4078 vdd.t106 vss 0.17868f
C4079 vdd.t107 vss 0.02206f
C4080 vdd.t214 vss 0.33339f
C4081 vdd.t360 vss 0.14187f
C4082 vdd.t305 vss 0.14187f
C4083 vdd.t326 vss 0.14187f
C4084 vdd.t327 vss 0.14187f
C4085 vdd.t367 vss 0.14187f
C4086 vdd.t223 vss 0.14187f
C4087 vdd.t213 vss 0.14187f
C4088 vdd.t276 vss 0.14187f
C4089 vdd.t318 vss 0.14187f
C4090 vdd.t422 vss 0.14187f
C4091 vdd.t354 vss 0.14187f
C4092 vdd.t319 vss 0.14187f
C4093 vdd.t359 vss 0.14187f
C4094 vdd.t355 vss 0.14187f
C4095 vdd.t277 vss 0.14187f
C4096 vdd.t224 vss 0.19365f
C4097 vdd.n207 vss 1.75279f
C4098 vdd.n208 vss 0.37876f
C4099 vdd.n209 vss 0.97858f
C4100 vdd.n210 vss 0.68724f
C4101 vdd.n211 vss 0.37876f
C4102 vdd.n212 vss 0.97858f
C4103 vdd.n213 vss 0.68724f
C4104 vdd.n214 vss 0.37876f
C4105 vdd.n215 vss 0.97858f
C4106 vdd.n216 vss 0.68724f
C4107 vdd.n217 vss 0.37876f
C4108 vdd.n218 vss 0.97858f
C4109 vdd.n219 vss 0.68724f
C4110 vdd.n220 vss 0.37876f
C4111 vdd.n221 vss 0.97858f
C4112 vdd.n222 vss 0.68724f
C4113 vdd.n223 vss 0.37876f
C4114 vdd.n224 vss 0.97858f
C4115 vdd.n225 vss 0.68724f
C4116 vdd.n226 vss 0.37876f
C4117 vdd.n227 vss 0.97858f
C4118 vdd.n228 vss 0.68724f
C4119 vdd.n229 vss 0.37876f
C4120 vdd.n230 vss 0.97858f
C4121 vdd.n231 vss 0.68724f
C4122 vdd.n232 vss 0.37876f
C4123 vdd.n233 vss 0.99052f
C4124 vdd.n234 vss 0.68724f
C4125 vdd.n235 vss 0.37876f
C4126 vdd.n236 vss 0.20093f
C4127 BUS[5].t22 vss 0.08272f
C4128 BUS[5].t17 vss 0.08272f
C4129 BUS[5].n0 vss 0.44552f
C4130 BUS[5].t19 vss 0.08272f
C4131 BUS[5].t21 vss 0.08272f
C4132 BUS[5].n1 vss 0.44289f
C4133 BUS[5].n2 vss 0.25937f
C4134 BUS[5].t20 vss 0.08272f
C4135 BUS[5].t18 vss 0.08272f
C4136 BUS[5].n3 vss 0.44289f
C4137 BUS[5].n4 vss 0.21881f
C4138 BUS[5].t11 vss 0.66732f
C4139 BUS[5].n5 vss 0.21139f
C4140 BUS[5].t4 vss 0.08272f
C4141 BUS[5].t7 vss 0.08272f
C4142 BUS[5].n6 vss 0.44813f
C4143 BUS[5].t14 vss 0.08272f
C4144 BUS[5].t16 vss 0.08272f
C4145 BUS[5].n7 vss 0.44556f
C4146 BUS[5].n8 vss 0.25349f
C4147 BUS[5].t8 vss 0.08272f
C4148 BUS[5].t15 vss 0.08272f
C4149 BUS[5].n9 vss 0.44556f
C4150 BUS[5].n10 vss 0.14712f
C4151 BUS[5].t0 vss 0.08272f
C4152 BUS[5].t2 vss 0.08272f
C4153 BUS[5].n11 vss 0.44556f
C4154 BUS[5].n12 vss 0.14712f
C4155 BUS[5].t5 vss 0.08272f
C4156 BUS[5].t12 vss 0.08272f
C4157 BUS[5].n13 vss 0.44556f
C4158 BUS[5].n14 vss 0.14712f
C4159 BUS[5].t3 vss 0.08272f
C4160 BUS[5].t6 vss 0.08272f
C4161 BUS[5].n15 vss 0.44556f
C4162 BUS[5].n16 vss 0.14712f
C4163 BUS[5].t13 vss 0.08272f
C4164 BUS[5].t10 vss 0.08272f
C4165 BUS[5].n17 vss 0.44556f
C4166 BUS[5].n18 vss 0.14712f
C4167 BUS[5].t1 vss 0.08272f
C4168 BUS[5].t9 vss 0.08272f
C4169 BUS[5].n19 vss 0.44556f
C4170 BUS[5].n20 vss 0.11197f
C4171 BUS[5].n21 vss 0.37951f
C4172 pin.t198 vss 0.5312f
C4173 pin.t195 vss 0.07503f
C4174 pin.t197 vss 0.07503f
C4175 pin.n0 vss 0.35364f
C4176 pin.t196 vss 0.07503f
C4177 pin.t199 vss 0.07503f
C4178 pin.n1 vss 0.35364f
C4179 pin.t194 vss 0.5312f
C4180 pin.t87 vss 0.07503f
C4181 pin.t228 vss 0.07503f
C4182 pin.n2 vss 0.35669f
C4183 pin.t118 vss 0.07503f
C4184 pin.t226 vss 0.07503f
C4185 pin.n3 vss 0.35669f
C4186 pin.t85 vss 0.07503f
C4187 pin.t50 vss 0.07503f
C4188 pin.n4 vss 0.35669f
C4189 pin.t51 vss 0.07503f
C4190 pin.t224 vss 0.07503f
C4191 pin.n5 vss 0.35669f
C4192 pin.t225 vss 0.07503f
C4193 pin.t86 vss 0.07503f
C4194 pin.n6 vss 0.35669f
C4195 pin.t119 vss 0.07503f
C4196 pin.t227 vss 0.07503f
C4197 pin.n7 vss 0.35669f
C4198 pin.t17 vss 0.07503f
C4199 pin.t16 vss 0.07503f
C4200 pin.n8 vss 0.35669f
C4201 pin.t88 vss 0.07503f
C4202 pin.t120 vss 0.07503f
C4203 pin.n9 vss 0.35669f
C4204 pin.t18 vss 0.5518f
C4205 pin.t68 vss 0.5312f
C4206 pin.t67 vss 0.07503f
C4207 pin.t65 vss 0.07503f
C4208 pin.n10 vss 0.35364f
C4209 pin.t64 vss 0.07503f
C4210 pin.t66 vss 0.07503f
C4211 pin.n11 vss 0.35364f
C4212 pin.t69 vss 0.5312f
C4213 pin.t5 vss 0.07503f
C4214 pin.t2 vss 0.07503f
C4215 pin.n12 vss 0.35669f
C4216 pin.t75 vss 0.07503f
C4217 pin.t43 vss 0.07503f
C4218 pin.n13 vss 0.35669f
C4219 pin.t8 vss 0.07503f
C4220 pin.t0 vss 0.07503f
C4221 pin.n14 vss 0.35669f
C4222 pin.t1 vss 0.07503f
C4223 pin.t76 vss 0.07503f
C4224 pin.n15 vss 0.35669f
C4225 pin.t57 vss 0.07503f
C4226 pin.t4 vss 0.07503f
C4227 pin.n16 vss 0.35669f
C4228 pin.t220 vss 0.07503f
C4229 pin.t82 vss 0.07503f
C4230 pin.n17 vss 0.35669f
C4231 pin.t9 vss 0.07503f
C4232 pin.t42 vss 0.07503f
C4233 pin.n18 vss 0.35669f
C4234 pin.t3 vss 0.07503f
C4235 pin.t77 vss 0.07503f
C4236 pin.n19 vss 0.35669f
C4237 pin.t56 vss 0.5518f
C4238 pin.t173 vss 0.5312f
C4239 pin.t174 vss 0.07503f
C4240 pin.t169 vss 0.07503f
C4241 pin.n20 vss 0.35364f
C4242 pin.t171 vss 0.07503f
C4243 pin.t172 vss 0.07503f
C4244 pin.n21 vss 0.35364f
C4245 pin.t170 vss 0.5312f
C4246 pin.t89 vss 0.07503f
C4247 pin.t53 vss 0.07503f
C4248 pin.n22 vss 0.35669f
C4249 pin.t95 vss 0.07503f
C4250 pin.t190 vss 0.07503f
C4251 pin.n23 vss 0.35669f
C4252 pin.t191 vss 0.07503f
C4253 pin.t52 vss 0.07503f
C4254 pin.n24 vss 0.35669f
C4255 pin.t93 vss 0.07503f
C4256 pin.t71 vss 0.07503f
C4257 pin.n25 vss 0.35669f
C4258 pin.t90 vss 0.07503f
C4259 pin.t20 vss 0.07503f
C4260 pin.n26 vss 0.35669f
C4261 pin.t21 vss 0.07503f
C4262 pin.t94 vss 0.07503f
C4263 pin.n27 vss 0.35669f
C4264 pin.t101 vss 0.07503f
C4265 pin.t91 vss 0.07503f
C4266 pin.n28 vss 0.35669f
C4267 pin.t19 vss 0.07503f
C4268 pin.t103 vss 0.07503f
C4269 pin.n29 vss 0.35669f
C4270 pin.t102 vss 0.5518f
C4271 pin.t202 vss 0.5312f
C4272 pin.t205 vss 0.07503f
C4273 pin.t201 vss 0.07503f
C4274 pin.n30 vss 0.35364f
C4275 pin.t200 vss 0.07503f
C4276 pin.t203 vss 0.07503f
C4277 pin.n31 vss 0.35364f
C4278 pin.t204 vss 0.5312f
C4279 pin.t128 vss 0.07503f
C4280 pin.t142 vss 0.07503f
C4281 pin.n32 vss 0.35669f
C4282 pin.t143 vss 0.07503f
C4283 pin.t107 vss 0.07503f
C4284 pin.n33 vss 0.35669f
C4285 pin.t132 vss 0.07503f
C4286 pin.t129 vss 0.07503f
C4287 pin.n34 vss 0.35669f
C4288 pin.t131 vss 0.07503f
C4289 pin.t168 vss 0.07503f
C4290 pin.n35 vss 0.35669f
C4291 pin.t141 vss 0.07503f
C4292 pin.t192 vss 0.07503f
C4293 pin.n36 vss 0.35669f
C4294 pin.t193 vss 0.07503f
C4295 pin.t159 vss 0.07503f
C4296 pin.n37 vss 0.35669f
C4297 pin.t133 vss 0.07503f
C4298 pin.t70 vss 0.07503f
C4299 pin.n38 vss 0.35669f
C4300 pin.t140 vss 0.07503f
C4301 pin.t130 vss 0.07503f
C4302 pin.n39 vss 0.35669f
C4303 pin.t167 vss 0.5518f
C4304 pin.t63 vss 0.5312f
C4305 pin.t59 vss 0.07503f
C4306 pin.t60 vss 0.07503f
C4307 pin.n40 vss 0.35364f
C4308 pin.t62 vss 0.07503f
C4309 pin.t58 vss 0.07503f
C4310 pin.n41 vss 0.35364f
C4311 pin.t61 vss 0.5312f
C4312 pin.t38 vss 0.07503f
C4313 pin.t35 vss 0.07503f
C4314 pin.n42 vss 0.35669f
C4315 pin.t34 vss 0.07503f
C4316 pin.t28 vss 0.07503f
C4317 pin.n43 vss 0.35669f
C4318 pin.t30 vss 0.07503f
C4319 pin.t26 vss 0.07503f
C4320 pin.n44 vss 0.35669f
C4321 pin.t40 vss 0.07503f
C4322 pin.t41 vss 0.07503f
C4323 pin.n45 vss 0.35669f
C4324 pin.t29 vss 0.07503f
C4325 pin.t33 vss 0.07503f
C4326 pin.n46 vss 0.35669f
C4327 pin.t31 vss 0.07503f
C4328 pin.t39 vss 0.07503f
C4329 pin.n47 vss 0.35669f
C4330 pin.t25 vss 0.07503f
C4331 pin.t37 vss 0.07503f
C4332 pin.n48 vss 0.35669f
C4333 pin.t32 vss 0.07503f
C4334 pin.t27 vss 0.07503f
C4335 pin.n49 vss 0.35669f
C4336 pin.t36 vss 0.5518f
C4337 pin.t176 vss 0.5312f
C4338 pin.t177 vss 0.07503f
C4339 pin.t180 vss 0.07503f
C4340 pin.n50 vss 0.35364f
C4341 pin.t179 vss 0.07503f
C4342 pin.t175 vss 0.07503f
C4343 pin.n51 vss 0.35364f
C4344 pin.t178 vss 0.5312f
C4345 pin.t117 vss 0.07503f
C4346 pin.t97 vss 0.07503f
C4347 pin.n52 vss 0.35669f
C4348 pin.t23 vss 0.07503f
C4349 pin.t153 vss 0.07503f
C4350 pin.n53 vss 0.35669f
C4351 pin.t183 vss 0.07503f
C4352 pin.t181 vss 0.07503f
C4353 pin.n54 vss 0.35669f
C4354 pin.t96 vss 0.07503f
C4355 pin.t24 vss 0.07503f
C4356 pin.n55 vss 0.35669f
C4357 pin.t152 vss 0.07503f
C4358 pin.t116 vss 0.07503f
C4359 pin.n56 vss 0.35669f
C4360 pin.t99 vss 0.07503f
C4361 pin.t154 vss 0.07503f
C4362 pin.n57 vss 0.35669f
C4363 pin.t22 vss 0.07503f
C4364 pin.t182 vss 0.07503f
C4365 pin.n58 vss 0.35669f
C4366 pin.t98 vss 0.07503f
C4367 pin.t100 vss 0.07503f
C4368 pin.n59 vss 0.35669f
C4369 pin.t212 vss 0.5518f
C4370 pin.t217 vss 0.5312f
C4371 pin.t218 vss 0.07503f
C4372 pin.t215 vss 0.07503f
C4373 pin.n60 vss 0.35364f
C4374 pin.t214 vss 0.07503f
C4375 pin.t216 vss 0.07503f
C4376 pin.n61 vss 0.35364f
C4377 pin.t213 vss 0.5312f
C4378 pin.t123 vss 0.07503f
C4379 pin.t145 vss 0.07503f
C4380 pin.n62 vss 0.35669f
C4381 pin.t222 vss 0.07503f
C4382 pin.t109 vss 0.07503f
C4383 pin.n63 vss 0.35669f
C4384 pin.t110 vss 0.07503f
C4385 pin.t219 vss 0.07503f
C4386 pin.n64 vss 0.35669f
C4387 pin.t149 vss 0.07503f
C4388 pin.t223 vss 0.07503f
C4389 pin.n65 vss 0.35669f
C4390 pin.t136 vss 0.07503f
C4391 pin.t151 vss 0.07503f
C4392 pin.n66 vss 0.35669f
C4393 pin.t122 vss 0.07503f
C4394 pin.t150 vss 0.07503f
C4395 pin.n67 vss 0.35669f
C4396 pin.t92 vss 0.07503f
C4397 pin.t137 vss 0.07503f
C4398 pin.n68 vss 0.35669f
C4399 pin.t165 vss 0.07503f
C4400 pin.t144 vss 0.07503f
C4401 pin.n69 vss 0.35669f
C4402 pin.t126 vss 0.5518f
C4403 pin.t13 vss 0.5312f
C4404 pin.t15 vss 0.07503f
C4405 pin.t10 vss 0.07503f
C4406 pin.n70 vss 0.35364f
C4407 pin.t12 vss 0.07503f
C4408 pin.t14 vss 0.07503f
C4409 pin.n71 vss 0.35364f
C4410 pin.t11 vss 0.5312f
C4411 pin.t114 vss 0.07503f
C4412 pin.t72 vss 0.07503f
C4413 pin.n72 vss 0.35669f
C4414 pin.t73 vss 0.07503f
C4415 pin.t104 vss 0.07503f
C4416 pin.n73 vss 0.35669f
C4417 pin.t105 vss 0.07503f
C4418 pin.t74 vss 0.07503f
C4419 pin.n74 vss 0.35669f
C4420 pin.t185 vss 0.07503f
C4421 pin.t55 vss 0.07503f
C4422 pin.n75 vss 0.35669f
C4423 pin.t115 vss 0.07503f
C4424 pin.t7 vss 0.07503f
C4425 pin.n76 vss 0.35669f
C4426 pin.t113 vss 0.07503f
C4427 pin.t186 vss 0.07503f
C4428 pin.n77 vss 0.35669f
C4429 pin.t106 vss 0.07503f
C4430 pin.t229 vss 0.07503f
C4431 pin.n78 vss 0.35669f
C4432 pin.t6 vss 0.07503f
C4433 pin.t184 vss 0.07503f
C4434 pin.n79 vss 0.35669f
C4435 pin.t54 vss 0.5518f
C4436 pin.t206 vss 0.5312f
C4437 pin.t208 vss 0.07503f
C4438 pin.t209 vss 0.07503f
C4439 pin.n80 vss 0.35364f
C4440 pin.t207 vss 0.07503f
C4441 pin.t210 vss 0.07503f
C4442 pin.n81 vss 0.35364f
C4443 pin.t211 vss 0.5312f
C4444 pin.t188 vss 0.07503f
C4445 pin.t135 vss 0.07503f
C4446 pin.n82 vss 0.35669f
C4447 pin.t108 vss 0.07503f
C4448 pin.t164 vss 0.07503f
C4449 pin.n83 vss 0.35669f
C4450 pin.t79 vss 0.07503f
C4451 pin.t125 vss 0.07503f
C4452 pin.n84 vss 0.35669f
C4453 pin.t221 vss 0.07503f
C4454 pin.t155 vss 0.07503f
C4455 pin.n85 vss 0.35669f
C4456 pin.t156 vss 0.07503f
C4457 pin.t187 vss 0.07503f
C4458 pin.n86 vss 0.35669f
C4459 pin.t148 vss 0.07503f
C4460 pin.t134 vss 0.07503f
C4461 pin.n87 vss 0.35669f
C4462 pin.t160 vss 0.07503f
C4463 pin.t121 vss 0.07503f
C4464 pin.n88 vss 0.35669f
C4465 pin.t78 vss 0.07503f
C4466 pin.t124 vss 0.07503f
C4467 pin.n89 vss 0.35669f
C4468 pin.t161 vss 0.5518f
C4469 pin.t49 vss 0.5312f
C4470 pin.t45 vss 0.07503f
C4471 pin.t46 vss 0.07503f
C4472 pin.n90 vss 0.35364f
C4473 pin.t47 vss 0.07503f
C4474 pin.t48 vss 0.07503f
C4475 pin.n91 vss 0.35364f
C4476 pin.t44 vss 0.5312f
C4477 pin.t163 vss 0.07503f
C4478 pin.t81 vss 0.07503f
C4479 pin.n92 vss 0.35669f
C4480 pin.t146 vss 0.07503f
C4481 pin.t127 vss 0.07503f
C4482 pin.n93 vss 0.35669f
C4483 pin.t166 vss 0.07503f
C4484 pin.t147 vss 0.07503f
C4485 pin.n94 vss 0.35669f
C4486 pin.t80 vss 0.07503f
C4487 pin.t83 vss 0.07503f
C4488 pin.n95 vss 0.35669f
C4489 pin.t138 vss 0.07503f
C4490 pin.t111 vss 0.07503f
C4491 pin.n96 vss 0.35669f
C4492 pin.t157 vss 0.07503f
C4493 pin.t189 vss 0.07503f
C4494 pin.n97 vss 0.35669f
C4495 pin.t162 vss 0.07503f
C4496 pin.t139 vss 0.07503f
C4497 pin.n98 vss 0.35669f
C4498 pin.t112 vss 0.07503f
C4499 pin.t158 vss 0.07503f
C4500 pin.n99 vss 0.35669f
C4501 pin.t84 vss 0.5667f
C4502 pin.n100 vss 1.02941f
C4503 pin.n101 vss 0.29021f
C4504 pin.n102 vss 0.29021f
C4505 pin.n103 vss 0.29021f
C4506 pin.n104 vss 0.29021f
C4507 pin.n105 vss 0.29021f
C4508 pin.n106 vss 0.29021f
C4509 pin.n107 vss 0.3977f
C4510 pin.n108 vss 0.43207f
C4511 pin.n109 vss 0.30013f
C4512 pin.n110 vss 0.29939f
C4513 pin.n111 vss 0.45703f
C4514 pin.n112 vss 0.50082f
C4515 pin.n113 vss 0.29762f
C4516 pin.n114 vss 0.29021f
C4517 pin.n115 vss 0.29021f
C4518 pin.n116 vss 0.29021f
C4519 pin.n117 vss 0.29021f
C4520 pin.n118 vss 0.29021f
C4521 pin.n119 vss 0.29021f
C4522 pin.n120 vss 0.3977f
C4523 pin.n121 vss 0.43207f
C4524 pin.n122 vss 0.30013f
C4525 pin.n123 vss 0.29939f
C4526 pin.n124 vss 0.45703f
C4527 pin.n125 vss 0.50082f
C4528 pin.n126 vss 0.29762f
C4529 pin.n127 vss 0.29021f
C4530 pin.n128 vss 0.29021f
C4531 pin.n129 vss 0.29021f
C4532 pin.n130 vss 0.29021f
C4533 pin.n131 vss 0.29021f
C4534 pin.n132 vss 0.29021f
C4535 pin.n133 vss 0.3977f
C4536 pin.n134 vss 0.43207f
C4537 pin.n135 vss 0.30013f
C4538 pin.n136 vss 0.29939f
C4539 pin.n137 vss 0.45703f
C4540 pin.n138 vss 0.50082f
C4541 pin.n139 vss 0.29762f
C4542 pin.n140 vss 0.29021f
C4543 pin.n141 vss 0.29021f
C4544 pin.n142 vss 0.29021f
C4545 pin.n143 vss 0.29021f
C4546 pin.n144 vss 0.29021f
C4547 pin.n145 vss 0.29021f
C4548 pin.n146 vss 0.3977f
C4549 pin.n147 vss 0.43207f
C4550 pin.n148 vss 0.30013f
C4551 pin.n149 vss 0.29939f
C4552 pin.n150 vss 0.45703f
C4553 pin.n151 vss 0.50082f
C4554 pin.n152 vss 0.29762f
C4555 pin.n153 vss 0.29021f
C4556 pin.n154 vss 0.29021f
C4557 pin.n155 vss 0.29021f
C4558 pin.n156 vss 0.29021f
C4559 pin.n157 vss 0.29021f
C4560 pin.n158 vss 0.29021f
C4561 pin.n159 vss 0.3977f
C4562 pin.n160 vss 0.43207f
C4563 pin.n161 vss 0.30013f
C4564 pin.n162 vss 0.29939f
C4565 pin.n163 vss 0.45703f
C4566 pin.n164 vss 0.50082f
C4567 pin.n165 vss 0.29762f
C4568 pin.n166 vss 0.29021f
C4569 pin.n167 vss 0.29021f
C4570 pin.n168 vss 0.29021f
C4571 pin.n169 vss 0.29021f
C4572 pin.n170 vss 0.29021f
C4573 pin.n171 vss 0.29021f
C4574 pin.n172 vss 0.3977f
C4575 pin.n173 vss 0.43207f
C4576 pin.n174 vss 0.30013f
C4577 pin.n175 vss 0.29939f
C4578 pin.n176 vss 0.45703f
C4579 pin.n177 vss 0.50082f
C4580 pin.n178 vss 0.29762f
C4581 pin.n179 vss 0.29021f
C4582 pin.n180 vss 0.29021f
C4583 pin.n181 vss 0.29021f
C4584 pin.n182 vss 0.29021f
C4585 pin.n183 vss 0.29021f
C4586 pin.n184 vss 0.29021f
C4587 pin.n185 vss 0.3977f
C4588 pin.n186 vss 0.43207f
C4589 pin.n187 vss 0.30013f
C4590 pin.n188 vss 0.29939f
C4591 pin.n189 vss 0.45703f
C4592 pin.n190 vss 0.50082f
C4593 pin.n191 vss 0.29762f
C4594 pin.n192 vss 0.29021f
C4595 pin.n193 vss 0.29021f
C4596 pin.n194 vss 0.29021f
C4597 pin.n195 vss 0.29021f
C4598 pin.n196 vss 0.29021f
C4599 pin.n197 vss 0.29021f
C4600 pin.n198 vss 0.3977f
C4601 pin.n199 vss 0.43207f
C4602 pin.n200 vss 0.30013f
C4603 pin.n201 vss 0.29939f
C4604 pin.n202 vss 0.45703f
C4605 pin.n203 vss 0.50082f
C4606 pin.n204 vss 0.29762f
C4607 pin.n205 vss 0.29021f
C4608 pin.n206 vss 0.29021f
C4609 pin.n207 vss 0.29021f
C4610 pin.n208 vss 0.29021f
C4611 pin.n209 vss 0.29021f
C4612 pin.n210 vss 0.29021f
C4613 pin.n211 vss 0.3977f
C4614 pin.n212 vss 0.43207f
C4615 pin.n213 vss 0.30013f
C4616 pin.n214 vss 0.29939f
C4617 pin.n215 vss 0.45703f
C4618 pin.n216 vss 0.52356f
C4619 pin.n217 vss 0.29762f
C4620 pin.n218 vss 0.29021f
C4621 pin.n219 vss 0.29021f
C4622 pin.n220 vss 0.29021f
C4623 pin.n221 vss 0.29021f
C4624 pin.n222 vss 0.29021f
C4625 pin.n223 vss 0.29021f
C4626 pin.n224 vss 0.3977f
C4627 pin.n225 vss 0.43207f
C4628 pin.n226 vss 0.30013f
C4629 pin.n227 vss 0.29939f
C4630 pin.n228 vss 0.45703f
C4631 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 vss 0.06945f
C4632 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 vss 0.09589f
C4633 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 vss 0.12443f
C4634 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 vss 0.1242f
C4635 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 vss 0.1906f
C4636 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 vss 0.1242f
C4637 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 vss 0.10127f
C4638 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 vss 0.1242f
C4639 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 vss 0.10127f
C4640 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 vss 0.1242f
C4641 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 vss 0.10127f
C4642 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 vss 0.1242f
C4643 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 vss 0.10127f
C4644 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 vss 0.1242f
C4645 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 vss 0.10127f
C4646 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 vss 0.1242f
C4647 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 vss 0.10127f
C4648 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 vss 0.1242f
C4649 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 vss 0.10127f
C4650 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 vss 0.1242f
C4651 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 vss 0.10127f
C4652 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 vss 0.1242f
C4653 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 vss 0.10127f
C4654 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 vss 0.1242f
C4655 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 vss 0.10127f
C4656 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 vss 0.1242f
C4657 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 vss 0.10127f
C4658 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 vss 0.1242f
C4659 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 vss 0.10127f
C4660 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 vss 0.1242f
C4661 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 vss 0.10127f
C4662 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 vss 0.1242f
C4663 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 vss 0.10127f
C4664 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 vss 0.1242f
C4665 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 vss 0.52842f
C4666 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 vss 0.49145f
.ends

