* NGSPICE file created from ah_syn_lifcomp.ext - technology: gf180mcuD

.subckt pfet$16 a_150_0# a_38_n60# a_n92_0# w_n230_n138#
X0 a_150_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.286p pd=2.18u as=0.286p ps=2.18u w=0.44u l=0.56u
.ends

.subckt nfet$32 a_n84_n2# a_194_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_194_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.78u
.ends

.subckt pfet$17 a_38_n60# a_n92_0# a_318_0# w_n230_n138#
X0 a_318_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=1.4u
.ends

.subckt nfet$30 a_150_0# dw_n710_n726# a_n84_0# a_38_n132# w_n710_n726#
X0 a_150_0# a_38_n132# a_n84_0# w_n710_n726# nfet_03v3 ad=0.2684p pd=2.1u as=0.2684p ps=2.1u w=0.44u l=0.56u
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=6u c_length=5u
.ends

.subckt nfet$33 a_1158_0# a_n84_n2# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_1158_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=5.6u
.ends

.subckt nfet$31 a_n84_n2# a_374_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_374_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=1.68u
.ends

.subckt AH_neuron$1 vdd Current_in v_bias vout vss
Xpfet$16_0 vdd Current_in m2_381_1901# vdd pfet$16
Xnfet$32_0 vout vss nfet$33_0/dw_n710_n726# m2_381_1901# vss nfet$32
Xpfet$17_0 m2_381_1901# vout vdd vdd pfet$17
Xnfet$30_0 vss nfet$33_0/dw_n710_n726# m2_381_1901# Current_in vss nfet$30
Xcap_mim$3_0 Current_in vout cap_mim$3
Xnfet$33_0 m1_335_n170# Current_in nfet$33_0/dw_n710_n726# v_bias vss nfet$33
Xnfet$31_0 m1_335_n170# vss nfet$33_0/dw_n710_n726# vout vss nfet$31
.ends

.subckt pfet$21 a_28_n136# w_n232_n142# a_94_0# a_n92_n2#
X0 a_94_0# a_28_n136# a_n92_n2# w_n232_n142# pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
.ends

.subckt nfet$36 dw_n710_n652# a_30_260# a_n84_0# a_94_0# w_n710_n652#
X0 a_94_0# a_30_260# a_n84_0# w_n710_n652# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$34 dw_n710_n726# a_30_n132# a_n84_0# a_94_0# w_n710_n726#
X0 a_94_0# a_30_n132# a_n84_0# w_n710_n726# nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$19 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
.ends

.subckt pfet$20 a_28_144# w_n232_n142# a_94_0# a_n92_n2#
X0 a_94_0# a_28_144# a_n92_n2# w_n232_n142# pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
.ends

.subckt nfet$37 a_n84_n2# dw_n710_n652# a_94_0# a_30_144# w_n710_n652#
X0 a_94_0# a_30_144# a_n84_n2# w_n710_n652# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
.ends

.subckt nfet$35 a_n84_n2# dw_n710_n726# a_30_n132# a_94_0# w_n710_n726#
X0 a_94_0# a_30_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
.ends

.subckt pfet$18 a_28_620# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_620# a_n92_0# w_n230_n138# pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
.ends

.subckt synapse vi v_ctrl v_in ve vdd v_out vss
Xpfet$21_0 vi vdd vdd m1_44_2533# pfet$21
Xnfet$36_0 nfet$37_0/dw_n710_n652# m1_344_2455# m1_2266_n82# vss vss nfet$36
Xnfet$34_0 nfet$37_0/dw_n710_n652# v_ctrl v_out m1_2266_n82# vss nfet$34
Xpfet$19_0 m2_640_1617# m1_1750_2493# vdd vdd pfet$19
Xpfet$20_0 v_in vdd vdd m1_856_n14# pfet$20
Xpfet$20_1 m1_856_n14# vdd m1_44_2533# m1_344_2455# pfet$20
Xnfet$37_0 m2_640_1617# nfet$37_0/dw_n710_n652# m1_1434_n778# v_in vss nfet$37
Xpfet$20_2 m2_640_1617# vdd vdd m2_640_1617# pfet$20
Xnfet$35_0 m1_1434_n778# nfet$37_0/dw_n710_n652# ve vss vss nfet$35
Xnfet$35_1 m1_856_n14# nfet$37_0/dw_n710_n652# v_in vss vss nfet$35
Xnfet$35_2 m1_344_2455# nfet$37_0/dw_n710_n652# m1_344_2455# vss vss nfet$35
Xpfet$18_0 v_ctrl v_out m1_1750_2493# vdd pfet$18
.ends

.subckt AH_neuron vdd Current_in v_bias vout vss
Xpfet$16_0 vdd Current_in m2_381_1901# vdd pfet$16
Xnfet$32_0 vout vss nfet$33_0/dw_n710_n726# m2_381_1901# vss nfet$32
Xpfet$17_0 m2_381_1901# vout vdd vdd pfet$17
Xnfet$30_0 vss nfet$33_0/dw_n710_n726# m2_381_1901# Current_in vss nfet$30
Xcap_mim$3_0 Current_in vout cap_mim$3
Xnfet$33_0 m1_335_n170# Current_in nfet$33_0/dw_n710_n726# v_bias vss nfet$33
Xnfet$31_0 m1_335_n170# vss nfet$33_0/dw_n710_n726# vout vss nfet$31
.ends

.subckt nfet$22 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$12 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt switch out cntrl in vdd vss
Xnfet$22_0 vss cntrl m2_n331_n296# vss nfet$22
Xnfet$22_1 vss cntrl in out nfet$22
Xpfet$12_0 m2_n331_n296# cntrl vdd vdd pfet$12
Xpfet$12_1 in m2_n331_n296# out vdd pfet$12
.ends

.subckt nfet$20 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$21 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt pfet$11 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$19 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_1stage vdd vp vn vss vout
Xnfet$20_0 vss vn m3_n530_n14# vout nfet$20
Xnfet$20_1 vss vp m3_n530_n14# m3_n314_178# nfet$20
Xnfet$21_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$21
Xnfet$21_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$21
Xpfet$11_0 vdd vdd m3_n314_178# m3_n314_178# pfet$11
Xpfet$11_1 vdd vdd vout m3_n314_178# pfet$11
Xnfet$19_0 m3_n1200_n476# vss vdd vdd nfet$19
.ends

.subckt cap_mim$2 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt nfet$29 a_n256_n198# a_38_n60# a_n84_0# a_138_0#
X0 a_138_0# a_38_n60# a_n84_0# a_n256_n198# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt pfet$14 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$27 a_n256_n198# a_30_228# a_n84_0# a_94_0#
X0 a_94_0# a_30_228# a_n84_0# a_n256_n198# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$25 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$15 a_28_n136# a_n92_0# a_94_0# w_n352_n362#
X0 a_94_0# a_28_n136# a_n92_0# w_n352_n362# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
.ends

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt nfet$28 a_n256_n198# a_30_172# a_n84_0# a_94_0#
X0 a_94_0# a_30_172# a_n84_0# a_n256_n198# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt nfet$26 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$24 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_2stage vdd vp vn vss vout
Xpfet$14_0 vdd vdd m3_n314_178# m3_n314_178# pfet$14
Xpfet$14_1 vdd m3_210_178# vdd m3_n314_178# pfet$14
Xnfet$27_0 vss m3_n1200_n227# m3_n1200_n227# vss nfet$27
Xnfet$25_0 vss vp m3_210_178# m3_n530_n14# nfet$25
Xnfet$25_1 vss vn m3_n530_n14# m3_n314_178# nfet$25
Xpfet$15_0 m3_210_178# vdd vout vdd pfet$15
Xcap_mim$1_0 vout m3_210_178# cap_mim$1
Xnfet$28_0 vss m3_n1200_n227# vss vout nfet$28
Xnfet$26_0 vss m3_n1200_n227# vss m3_n530_n14# nfet$26
Xnfet$24_0 m3_n1200_n227# vss vdd vdd nfet$24
.ends

.subckt nfet$23 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$13 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt conmutator in1 in2 vdd out cntrl vss
Xnfet$23_0 vss m2_n850_n472# out in1 nfet$23
Xnfet$23_1 vss cntrl in2 out nfet$23
Xnfet$23_2 vss cntrl m2_n850_n472# vss nfet$23
Xpfet$13_0 out cntrl in1 vdd pfet$13
Xpfet$13_2 m2_n850_n472# cntrl vdd vdd pfet$13
Xpfet$13_1 in2 m2_n850_n472# out vdd pfet$13
.ends

.subckt nfet$9 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.3355p pd=2.32u as=0.3355p ps=2.32u w=0.55u l=0.28u
.ends

.subckt nfet$7 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$8 a_n256_n272# a_n84_0# a_198_0# a_38_n132#
X0 a_198_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.8u
.ends

.subckt nfet$6 a_n84_n2# a_n256_n272# a_30_n132# a_94_0#
X0 a_94_0# a_30_n132# a_n84_n2# a_n256_n272# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
.ends

.subckt nvdiv vss vdd vspike_up vspike_down vres vref
Xnfet$9_0 vss vdd vdd vref nfet$9
Xnfet$7_0 vss vspike_down vspike_down vres nfet$7
Xnfet$7_1 vss m2_367_1540# m2_367_1540# vspike_down nfet$7
Xnfet$8_0 vss vres vss vres nfet$8
Xnfet$6_0 vref vss vref vss nfet$6
Xnfet$6_1 vspike_up vss vspike_up m2_367_1540# nfet$6
Xnfet$6_2 vdd vss vdd vspike_up nfet$6
.ends

.subckt pfet$7 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$12 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt not$1 out in vdd vss
Xpfet$7_0 out in vdd vdd pfet$7
Xnfet$12_0 vss in out vss nfet$12
.ends

.subckt pfet$6 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$11 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt switch$1 cntrl in vdd vss out
Xpfet$6_0 m2_n331_n296# cntrl vdd vdd pfet$6
Xpfet$6_1 in m2_n331_n296# out vdd pfet$6
Xnfet$11_0 vss cntrl m2_n331_n296# vss nfet$11
Xnfet$11_1 vss cntrl in out nfet$11
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt nfet$18 a_98_0# a_n256_n272# a_n84_0# a_32_n132#
X0 a_98_0# a_32_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
.ends

.subckt nfet$3 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$1 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt not out in vdd vss
Xnfet$3_0 vss in out vss nfet$3
Xpfet$1_0 out in vdd vdd pfet$1
.ends

.subckt pfet$4 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$5 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$3 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$4 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nand A B Z vdd vss
Xpfet$4_0 B Z vdd vdd pfet$4
Xnfet$5_0 A Z nfet$5_0/a_94_0# vss nfet$5
Xpfet$3_0 A vdd vdd Z pfet$3
Xnfet$4_0 vss B nfet$5_0/a_94_0# vss nfet$4
.ends

.subckt monostable vin vres phi_1 vneg vdd vss phi_2
Xcap_mim_0 not_1/in nand_0/Z cap_mim
Xcap_mim_1 not_3/in nand_1/Z cap_mim
Xnfet$18_0 vss vss not_1/in vres nfet$18
Xnot_0 phi_2 not_0/in vdd vss not
Xnfet$18_1 vss vss not_3/in vres nfet$18
Xnot_1 not_0/in not_1/in vdd vss not
Xnot_2 phi_1 vneg vdd vss not
Xnot_3 vneg not_3/in vdd vss not
Xnand_0 not_0/in phi_1 nand_0/Z vdd vss nand
Xnand_1 vneg vin nand_1/Z vdd vss nand
.ends

.subckt nfet$13 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$10 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt pfet$9 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$14 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nor A B Z vdd vss
Xnfet$13_0 vss A Z vss nfet$13
Xpfet$10_0 A pfet$9_0/a_94_0# vdd vdd pfet$10
Xpfet$9_0 B vdd Z pfet$9_0/a_94_0# pfet$9
Xnfet$14_0 B vss Z vss nfet$14
.ends

.subckt pfet$5 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$10 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$1 out in1 in2 vdd cntrl vss
Xpfet$5_0 out cntrl in1 vdd pfet$5
Xpfet$5_1 in2 m2_n850_n472# out vdd pfet$5
Xpfet$5_2 m2_n850_n472# cntrl vdd vdd pfet$5
Xnfet$10_0 vss m2_n850_n472# out in1 nfet$10
Xnfet$10_1 vss cntrl in2 out nfet$10
Xnfet$10_2 vss cntrl m2_n850_n472# vss nfet$10
.ends

.subckt nfet$17 a_2638_0# a_n84_n2# a_n256_n198# a_38_n60#
X0 a_2638_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=13u
.ends

.subckt nfet$15 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$16 a_n256_n198# a_30_3060# a_n84_0# a_94_0#
X0 a_94_0# a_30_3060# a_n84_0# a_n256_n198# nfet_03v3 ad=9.15p pd=31.22u as=9.15p ps=31.22u w=15u l=0.28u
.ends

.subckt pfet w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$1 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt nfet$2 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt ota_1stage$1 vdd vp vn vss vout
Xpfet_0 vdd vdd m3_n314_178# m3_n314_178# pfet
Xpfet_1 vdd vdd vout m3_n314_178# pfet
Xnfet$1_0 vss vn m3_n530_n14# vout nfet$1
Xnfet$1_1 vss vp m3_n530_n14# m3_n314_178# nfet$1
Xnfet_0 m3_n1200_n476# vss vdd vdd nfet
Xnfet$2_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$2
Xnfet$2_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$2
.ends

.subckt refractory vneg vss vspike_down vdd vrefrac
Xnfet$17_0 vneg ota_1stage$1_0/vp vss vneg nfet$17
Xnfet$15_0 vss ota_1stage$1_0/vn vspike_down vspike_down nfet$15
Xnfet$15_1 vss ota_1stage$1_0/vn ota_1stage$1_0/vn vrefrac nfet$15
Xnfet$16_0 vss ota_1stage$1_0/vp vss ota_1stage$1_0/vp nfet$16
Xota_1stage$1_0 vdd ota_1stage$1_0/vp ota_1stage$1_0/vn vss vrefrac ota_1stage$1
.ends

.subckt phaseUpulse phi_fire vin vspike reward vres vdd vref vss
Xnvdiv_0 vss vdd vspike_up vspike_down vres vref nvdiv
Xnot$1_0 phi_fire phi_int vdd vss not$1
Xswitch$1_0 phi_1 vspike vdd vss switch$1_0/out switch$1
Xswitch$1_1 phi_2 vspike vdd vss vrefrac switch$1
Xmonostable_0 vin vres phi_1 vneg vdd vss phi_2 monostable
Xswitch$1_2 phi_int vspike vdd vss vref switch$1
Xnor_0 phi_1 phi_2 phi_int vdd vss nor
Xconmutator$1_0 switch$1_0/out vspike_up vdd vdd reward vss conmutator$1
Xrefractory_0 vneg vss vspike_down vdd vrefrac refractory
.ends

.subckt LIF_comp vdd vin v_rew vout vss
Xswitch_0 vmem phi_fire vin vdd vss switch
Xota_1stage_0 vdd ota_1stage_0/vp v_th vss phaseUpulse_0/vin ota_1stage
Xcap_mim$2_0 conmutator_2/out vin cap_mim$2
Xnfet$29_0 vss v_th vin vmem nfet$29
Xota_2stage_0 vdd vspike vin vss vmem ota_2stage
Xconmutator_0 vmem vss vdd ota_1stage_0/vp phi_fire vss conmutator
Xconmutator_1 v_ref vmem vdd vout phi_fire vss conmutator
Xconmutator_2 vmem v_ref vdd conmutator_2/out phi_fire vss conmutator
XphaseUpulse_0 phi_fire phaseUpulse_0/vin vspike v_rew v_th vdd v_ref vss phaseUpulse
.ends

.subckt ah_syn_lifcomp vss vdd vout_lif vin_lif i_in0 vout_0 i_in1 vout_1 i_in2 vout_2
+ i_in3 vout_3 i_in4 vout_4 VAH_bias v_ex v_inh vin_s0 vout_s0 vin_s1 vout_s1 vin_s2
+ vout_s2 vin_s3 vout_s3 vin_s4 vout_s4 vin_s5 vout_s5
XAH_neuron$1_0 vdd i_in1 VAH_bias vout_1 vss AH_neuron$1
XAH_neuron$1_1 vdd i_in3 VAH_bias vout_3 vss AH_neuron$1
XAH_neuron$1_2 vdd i_in2 VAH_bias vout_2 vss AH_neuron$1
XAH_neuron$1_3 vdd i_in0 VAH_bias vout_0 vss AH_neuron$1
Xsynapse_0 v_inh synapse_0/v_ctrl vin_s1 v_ex vdd vout_s1 vss synapse
Xsynapse_1 v_inh synapse_1/v_ctrl vin_s0 v_ex vdd vout_s0 vss synapse
Xsynapse_2 v_inh synapse_2/v_ctrl vin_s4 v_ex vdd vout_s4 vss synapse
Xsynapse_3 v_inh synapse_3/v_ctrl vin_s5 v_ex vdd vout_s5 vss synapse
XAH_neuron_0 vdd i_in4 VAH_bias vout_4 vss AH_neuron
XLIF_comp_0 vdd vin_lif vss vout_lif vss LIF_comp
Xsynapse_4 v_inh synapse_4/v_ctrl vin_s2 v_ex vdd vout_s2 vss synapse
Xsynapse_5 v_inh synapse_5/v_ctrl vin_s3 v_ex vdd vout_s3 vss synapse
.ends

