* NGSPICE file created from swmatrix_Tgate.ext - technology: gf180mcuD
.subckt swmatrix_Tgate_pex gated_control T2 T1 VSS VDD
X0 VDD.t1 gated_control.t0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 VDD.t0 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 T1.t23 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 T2.t6 VDD.t19 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X2 T2.t9 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 T1.t22 VDD.t18 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X3 T2.t15 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 T1.t21 VDD.t17 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X4 T1.t20 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 T2.t18 VDD.t16 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X5 T1.t5 gated_control.t1 T2.t1 VSS.t7 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X6 T2.t3 gated_control.t2 T1.t4 VSS.t6 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X7 T1.t19 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 T2.t19 VDD.t15 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X8 T1.t18 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 T2.t21 VDD.t14 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X9 T2.t10 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 T1.t17 VDD.t13 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X10 T1.t16 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 T2.t16 VDD.t12 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X11 T2.t4 gated_control.t3 T1.t3 VSS.t5 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X12 T1.t2 gated_control.t4 T2.t5 VSS.t4 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X13 T2.t23 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 T1.t15 VDD.t11 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X14 T2.t22 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 T1.t14 VDD.t10 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X15 VSS.t3 gated_control.t5 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 VSS.t2 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X16 T2.t20 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 T1.t13 VDD.t9 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X17 T1.t12 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 T2.t13 VDD.t8 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X18 T2.t7 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 T1.t11 VDD.t7 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X19 T1.t10 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 T2.t11 VDD.t6 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X20 T2.t0 gated_control.t6 T1.t1 VSS.t1 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X21 T2.t17 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 T1.t9 VDD.t5 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X22 T1.t0 gated_control.t7 T2.t2 VSS.t0 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X23 T1.t8 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 T2.t14 VDD.t4 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X24 T2.t8 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 T1.t7 VDD.t3 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X25 T1.t6 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t19 T2.t12 VDD.t2 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
R0 gated_control.n1 gated_control.t4 71.7971
R1 gated_control.n5 gated_control.t6 71.6148
R2 gated_control.n4 gated_control.t1 71.6148
R3 gated_control.n3 gated_control.t3 71.6148
R4 gated_control.n2 gated_control.t7 71.6148
R5 gated_control.n1 gated_control.t2 71.6148
R6 gated_control.n0 gated_control.t0 23.3605
R7 gated_control.n0 gated_control.t5 15.2818
R8 gated_control gated_control.n5 5.96029
R9 gated_control.n6 gated_control 4.91117
R10 gated_control.n6 gated_control.n0 4.0128
R11 gated_control.n2 gated_control.n1 0.182778
R12 gated_control.n3 gated_control.n2 0.182778
R13 gated_control.n4 gated_control.n3 0.182778
R14 gated_control.n5 gated_control.n4 0.182778
R15 gated_control gated_control.n6 0.016687
R16 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 71.7994
R17 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 71.6148
R18 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 71.6148
R19 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 71.6148
R20 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t19 71.6148
R21 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 71.6148
R22 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 71.6148
R23 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 71.6148
R24 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 71.6148
R25 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 71.6148
R26 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 71.6148
R27 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 71.6148
R28 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 71.6148
R29 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 71.6148
R30 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 71.6148
R31 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 71.6148
R32 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 71.6148
R33 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 71.6148
R34 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n17 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 11.4757
R35 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 4.63372
R36 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n17 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 3.85252
R37 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n17 0.402556
R38 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 0.185115
R39 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 0.185115
R40 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 0.185115
R41 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 0.185115
R42 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 0.185115
R43 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 0.185115
R44 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 0.185115
R45 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 0.185115
R46 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 0.185115
R47 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 0.185115
R48 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 0.185115
R49 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 0.185115
R50 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 0.185115
R51 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 0.185115
R52 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 0.185115
R53 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 0.185115
R54 VDD.n1 VDD.t0 652.42
R55 VDD.n0 VDD.t4 245.306
R56 VDD.t0 VDD 195.008
R57 VDD.t4 VDD.t11 148.7
R58 VDD.t11 VDD.t15 148.7
R59 VDD.t15 VDD.t18 148.7
R60 VDD.t18 VDD.t8 148.7
R61 VDD.t8 VDD.t10 148.7
R62 VDD.t10 VDD.t19 148.7
R63 VDD.t19 VDD.t9 148.7
R64 VDD.t9 VDD.t6 148.7
R65 VDD.t6 VDD.t13 148.7
R66 VDD.t13 VDD.t16 148.7
R67 VDD.t16 VDD.t7 148.7
R68 VDD.t7 VDD.t14 148.7
R69 VDD.t14 VDD.t17 148.7
R70 VDD.t17 VDD.t2 148.7
R71 VDD.t2 VDD.t5 148.7
R72 VDD.t5 VDD.t12 148.7
R73 VDD.t12 VDD.t3 148.7
R74 VDD.n0 VDD.t1 3.84351
R75 VDD VDD.n1 0.0919062
R76 VDD VDD.n0 0.037625
R77 VDD.n1 VDD 0.001625
R78 T2.n2 T2.n0 15.3751
R79 T2.n9 T2.n7 15.2168
R80 T2.n2 T2.n1 15.0151
R81 T2.n4 T2.n3 15.0151
R82 T2.n21 T2.n20 14.8568
R83 T2.n19 T2.n18 14.8568
R84 T2.n17 T2.n16 14.8568
R85 T2.n15 T2.n14 14.8568
R86 T2.n13 T2.n12 14.8568
R87 T2.n11 T2.n10 14.8568
R88 T2.n9 T2.n8 14.8568
R89 T2.n6 T2.n5 14.8568
R90 T2.n6 T2.n4 0.8825
R91 T2.n20 T2.t12 0.4555
R92 T2.n20 T2.t17 0.4555
R93 T2.n18 T2.t21 0.4555
R94 T2.n18 T2.t15 0.4555
R95 T2.n16 T2.t18 0.4555
R96 T2.n16 T2.t7 0.4555
R97 T2.n14 T2.t11 0.4555
R98 T2.n14 T2.t10 0.4555
R99 T2.n12 T2.t6 0.4555
R100 T2.n12 T2.t20 0.4555
R101 T2.n10 T2.t13 0.4555
R102 T2.n10 T2.t22 0.4555
R103 T2.n8 T2.t19 0.4555
R104 T2.n8 T2.t9 0.4555
R105 T2.n7 T2.t14 0.4555
R106 T2.n7 T2.t23 0.4555
R107 T2.n5 T2.t16 0.4555
R108 T2.n5 T2.t8 0.4555
R109 T2.n0 T2.t1 0.41
R110 T2.n0 T2.t0 0.41
R111 T2.n1 T2.t2 0.41
R112 T2.n1 T2.t4 0.41
R113 T2.n3 T2.t5 0.41
R114 T2.n3 T2.t3 0.41
R115 T2.n4 T2.n2 0.3605
R116 T2.n11 T2.n9 0.3605
R117 T2.n13 T2.n11 0.3605
R118 T2.n15 T2.n13 0.3605
R119 T2.n17 T2.n15 0.3605
R120 T2.n19 T2.n17 0.3605
R121 T2.n21 T2.n19 0.3605
R122 T2.n22 T2.n6 0.219875
R123 T2 T2.n22 0.0545
R124 T2.n22 T2.n21 0.028625
R125 T1.n10 T1.t8 11.6271
R126 T1.n19 T1.t2 11.3631
R127 T1.n22 T1.t1 11.3631
R128 T1.n18 T1.t7 11.3121
R129 T1.n20 T1.n1 10.7331
R130 T1.n21 T1.n0 10.7331
R131 T1.n10 T1.n9 10.5771
R132 T1.n11 T1.n8 10.5771
R133 T1.n12 T1.n7 10.5771
R134 T1.n13 T1.n6 10.5771
R135 T1.n14 T1.n5 10.5771
R136 T1.n15 T1.n4 10.5771
R137 T1.n16 T1.n3 10.5771
R138 T1.n17 T1.n2 10.5771
R139 T1 T1.n22 0.7736
R140 T1.n9 T1.t15 0.4555
R141 T1.n9 T1.t19 0.4555
R142 T1.n8 T1.t22 0.4555
R143 T1.n8 T1.t12 0.4555
R144 T1.n7 T1.t14 0.4555
R145 T1.n7 T1.t23 0.4555
R146 T1.n6 T1.t13 0.4555
R147 T1.n6 T1.t10 0.4555
R148 T1.n5 T1.t17 0.4555
R149 T1.n5 T1.t20 0.4555
R150 T1.n4 T1.t11 0.4555
R151 T1.n4 T1.t18 0.4555
R152 T1.n3 T1.t21 0.4555
R153 T1.n3 T1.t6 0.4555
R154 T1.n2 T1.t9 0.4555
R155 T1.n2 T1.t16 0.4555
R156 T1.n1 T1.t4 0.41
R157 T1.n1 T1.t0 0.41
R158 T1.n0 T1.t3 0.41
R159 T1.n0 T1.t5 0.41
R160 T1.n19 T1.n18 0.365
R161 T1.n18 T1.n17 0.3155
R162 T1.n20 T1.n19 0.3146
R163 T1.n22 T1.n21 0.3119
R164 T1.n11 T1.n10 0.2885
R165 T1.n12 T1.n11 0.2885
R166 T1.n13 T1.n12 0.2885
R167 T1.n14 T1.n13 0.2885
R168 T1.n15 T1.n14 0.2885
R169 T1.n16 T1.n15 0.2885
R170 T1.n17 T1.n16 0.2885
R171 T1.n21 T1.n20 0.2885
R172 VSS.n1 VSS.t2 2022.85
R173 VSS VSS.t1 1140.15
R174 VSS.t4 VSS 554.961
R175 VSS.t2 VSS 551.977
R176 VSS.t6 VSS.t4 354.224
R177 VSS.t0 VSS.t6 354.224
R178 VSS.t5 VSS.t0 354.224
R179 VSS.t7 VSS.t5 354.224
R180 VSS.t1 VSS.t7 354.224
R181 VSS.n0 VSS.t3 4.63989
R182 VSS VSS.n0 1.64352
R183 VSS VSS.n1 0.0632187
R184 VSS VSS.n0 0.04325
R185 VSS.n1 VSS 0.001625
C0 gated_control VDD 1.51813f
C1 gated_control gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 0.8363f
C2 T1 T2 10.9994f
C3 T2 VDD 0.43357f
C4 T1 VDD 0.97222f
C5 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN T2 1.22075f
C6 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN 1.5419f
C7 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN VDD 5.07517f
C8 gated_control T2 0.34844f
C9 a_5322_453# VDD 0.00618f
C10 T1 gated_control 0.60389f
C11 T2 VSS 2.9617f
C12 T1 VSS 2.82624f
C13 gated_control VSS 1.89479f
C14 VDD VSS 15.44543f
C15 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN VSS 1.92827f
C16 T1.t1 VSS 0.51997f
C17 T1.t3 VSS 0.0734f
C18 T1.t5 VSS 0.0734f
C19 T1.n0 VSS 0.34623f
C20 T1.t4 VSS 0.0734f
C21 T1.t0 VSS 0.0734f
C22 T1.n1 VSS 0.34623f
C23 T1.t2 VSS 0.51997f
C24 T1.t7 VSS 0.54013f
C25 T1.t9 VSS 0.0734f
C26 T1.t16 VSS 0.0734f
C27 T1.n2 VSS 0.34921f
C28 T1.t21 VSS 0.0734f
C29 T1.t6 VSS 0.0734f
C30 T1.n3 VSS 0.34921f
C31 T1.t11 VSS 0.0734f
C32 T1.t18 VSS 0.0734f
C33 T1.n4 VSS 0.34921f
C34 T1.t17 VSS 0.0734f
C35 T1.t20 VSS 0.0734f
C36 T1.n5 VSS 0.34921f
C37 T1.t13 VSS 0.0734f
C38 T1.t10 VSS 0.0734f
C39 T1.n6 VSS 0.34921f
C40 T1.t14 VSS 0.0734f
C41 T1.t23 VSS 0.0734f
C42 T1.n7 VSS 0.34921f
C43 T1.t22 VSS 0.0734f
C44 T1.t12 VSS 0.0734f
C45 T1.n8 VSS 0.34921f
C46 T1.t15 VSS 0.0734f
C47 T1.t19 VSS 0.0734f
C48 T1.n9 VSS 0.34921f
C49 T1.t8 VSS 0.54842f
C50 T1.n10 VSS 0.55004f
C51 T1.n11 VSS 0.24723f
C52 T1.n12 VSS 0.24723f
C53 T1.n13 VSS 0.24723f
C54 T1.n14 VSS 0.24723f
C55 T1.n15 VSS 0.24723f
C56 T1.n16 VSS 0.24723f
C57 T1.n17 VSS 0.25252f
C58 T1.n18 VSS 0.29681f
C59 T1.n19 VSS 0.29393f
C60 T1.n20 VSS 0.25504f
C61 T1.n21 VSS 0.25451f
C62 T1.n22 VSS 0.37351f
C63 T2.t1 VSS 0.10179f
C64 T2.t0 VSS 0.10179f
C65 T2.n0 VSS 0.54819f
C66 T2.t2 VSS 0.10179f
C67 T2.t4 VSS 0.10179f
C68 T2.n1 VSS 0.54496f
C69 T2.n2 VSS 0.31915f
C70 T2.t5 VSS 0.10179f
C71 T2.t3 VSS 0.10179f
C72 T2.n3 VSS 0.54496f
C73 T2.n4 VSS 0.2755f
C74 T2.t16 VSS 0.10179f
C75 T2.t8 VSS 0.10179f
C76 T2.n5 VSS 0.54824f
C77 T2.n6 VSS 0.24739f
C78 T2.t14 VSS 0.10179f
C79 T2.t23 VSS 0.10179f
C80 T2.n7 VSS 0.55141f
C81 T2.t19 VSS 0.10179f
C82 T2.t9 VSS 0.10179f
C83 T2.n8 VSS 0.54824f
C84 T2.n9 VSS 0.31191f
C85 T2.t13 VSS 0.10179f
C86 T2.t22 VSS 0.10179f
C87 T2.n10 VSS 0.54824f
C88 T2.n11 VSS 0.18103f
C89 T2.t6 VSS 0.10179f
C90 T2.t20 VSS 0.10179f
C91 T2.n12 VSS 0.54824f
C92 T2.n13 VSS 0.18103f
C93 T2.t11 VSS 0.10179f
C94 T2.t10 VSS 0.10179f
C95 T2.n14 VSS 0.54824f
C96 T2.n15 VSS 0.18103f
C97 T2.t18 VSS 0.10179f
C98 T2.t7 VSS 0.10179f
C99 T2.n16 VSS 0.54824f
C100 T2.n17 VSS 0.18103f
C101 T2.t21 VSS 0.10179f
C102 T2.t15 VSS 0.10179f
C103 T2.n18 VSS 0.54824f
C104 T2.n19 VSS 0.18103f
C105 T2.t12 VSS 0.10179f
C106 T2.t17 VSS 0.10179f
C107 T2.n20 VSS 0.54824f
C108 T2.n21 VSS 0.12329f
C109 T2.n22 VSS -0.29221f
C110 VDD.t1 VSS 0.02612f
C111 VDD.t3 VSS 0.39481f
C112 VDD.t12 VSS 0.16801f
C113 VDD.t5 VSS 0.16801f
C114 VDD.t2 VSS 0.16801f
C115 VDD.t17 VSS 0.16801f
C116 VDD.t14 VSS 0.16801f
C117 VDD.t7 VSS 0.16801f
C118 VDD.t16 VSS 0.16801f
C119 VDD.t13 VSS 0.16801f
C120 VDD.t6 VSS 0.16801f
C121 VDD.t9 VSS 0.16801f
C122 VDD.t19 VSS 0.16801f
C123 VDD.t10 VSS 0.16801f
C124 VDD.t8 VSS 0.16801f
C125 VDD.t18 VSS 0.16801f
C126 VDD.t15 VSS 0.16801f
C127 VDD.t11 VSS 0.16801f
C128 VDD.t4 VSS 0.22975f
C129 VDD.n0 VSS 0.98121f
C130 VDD.t0 VSS 0.1711f
C131 VDD.n1 VSS 0.34748f
C132 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t1 VSS 0.06869f
C133 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t0 VSS 0.09485f
C134 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t17 VSS 0.12308f
C135 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t10 VSS 0.12285f
C136 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n0 VSS 0.18852f
C137 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t6 VSS 0.12285f
C138 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n1 VSS 0.10017f
C139 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t3 VSS 0.12285f
C140 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n2 VSS 0.10017f
C141 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t13 VSS 0.12285f
C142 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n3 VSS 0.10017f
C143 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t11 VSS 0.12285f
C144 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n4 VSS 0.10017f
C145 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t2 VSS 0.12285f
C146 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n5 VSS 0.10017f
C147 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t12 VSS 0.12285f
C148 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n6 VSS 0.10017f
C149 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t15 VSS 0.12285f
C150 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n7 VSS 0.10017f
C151 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t8 VSS 0.12285f
C152 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n8 VSS 0.10017f
C153 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t5 VSS 0.12285f
C154 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n9 VSS 0.10017f
C155 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t14 VSS 0.12285f
C156 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n10 VSS 0.10017f
C157 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t7 VSS 0.12285f
C158 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n11 VSS 0.10017f
C159 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t4 VSS 0.12285f
C160 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n12 VSS 0.10017f
C161 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t19 VSS 0.12285f
C162 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n13 VSS 0.10017f
C163 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t16 VSS 0.12285f
C164 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n14 VSS 0.10017f
C165 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t9 VSS 0.12285f
C166 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n15 VSS 0.10017f
C167 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.t18 VSS 0.12285f
C168 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n16 VSS 0.47233f
C169 gf180mcu_fd_sc_mcu9t5v0__inv_1_0.ZN.n17 VSS 0.46794f
.ends

