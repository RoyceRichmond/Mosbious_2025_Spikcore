* NGSPICE file created from LIF_comp.ext - technology: gf180mcuD

<<<<<<< HEAD
.subckt pfet w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$1 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt nfet$2 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt ota_1stage$2 vdd vp vn vss vout
Xpfet_0 vdd vdd m3_n314_178# m3_n314_178# pfet
Xpfet_1 vdd vdd vout m3_n314_178# pfet
Xnfet$1_0 vss vn m3_n530_n14# vout nfet$1
Xnfet$1_1 vss vp m3_n530_n14# m3_n314_178# nfet$1
Xnfet_0 m3_n1200_n476# vss vdd vdd nfet
Xnfet$2_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$2
Xnfet$2_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$2
.ends

.subckt nfet$50 a_n256_n198# a_38_n60# a_n84_0# a_138_0#
X0 a_138_0# a_38_n60# a_n84_0# a_n256_n198# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt pfet$16 a_28_n136# a_n92_0# a_94_0# w_n352_n362#
X0 a_94_0# a_28_n136# a_n92_0# w_n352_n362# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
.ends

.subckt nfet$27 a_n256_n198# a_30_228# a_n84_0# a_94_0#
X0 a_94_0# a_30_228# a_n84_0# a_n256_n198# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$25 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$15 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt nfet$28 a_n256_n198# a_30_172# a_n84_0# a_94_0#
X0 a_94_0# a_30_172# a_n84_0# a_n256_n198# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt nfet$26 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$24 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_2stage vdd vp vn vss vout
Xpfet$16_0 m3_210_178# vdd vout vdd pfet$16
Xnfet$27_0 vss m3_n1200_n227# m3_n1200_n227# vss nfet$27
Xnfet$25_0 vss vp m3_210_178# m3_n530_n14# nfet$25
Xnfet$25_1 vss vn m3_n530_n14# m3_n314_178# nfet$25
Xpfet$15_0 vdd vdd m3_n314_178# m3_n314_178# pfet$15
Xpfet$15_1 vdd m3_210_178# vdd m3_n314_178# pfet$15
Xcap_mim$1_0 vout m3_210_178# cap_mim$1
Xnfet$28_0 vss m3_n1200_n227# vss vout nfet$28
Xnfet$26_0 vss m3_n1200_n227# vss m3_n530_n14# nfet$26
Xnfet$24_0 m3_n1200_n227# vss vdd vdd nfet$24
.ends

.subckt pfet$6 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$11 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt switch$1 out cntrl in vdd vss
Xpfet$6_0 m2_n331_n296# cntrl vdd vdd pfet$6
Xpfet$6_1 in m2_n331_n296# out vdd pfet$6
Xnfet$11_0 vss cntrl m2_n331_n296# vss nfet$11
Xnfet$11_1 vss cntrl in out nfet$11
.ends

.subckt pfet$5 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$10 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$1 in1 in2 vdd out cntrl vss
Xpfet$5_0 out cntrl in1 vdd pfet$5
Xpfet$5_1 in2 m2_n850_n472# out vdd pfet$5
Xpfet$5_2 m2_n850_n472# cntrl vdd vdd pfet$5
Xnfet$10_0 vss m2_n850_n472# out in1 nfet$10
Xnfet$10_1 vss cntrl in2 out nfet$10
Xnfet$10_2 vss cntrl m2_n850_n472# vss nfet$10
=======
.subckt cap_mim$4 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt ppolyf_u_resistor$3 a_n376_0# a_160_0# a_n132_0#
X0 a_n132_0# a_160_0# a_n376_0# ppolyf_u r_width=0.8u r_length=0.8u
.ends

.subckt vdiv$1 vss vspike_up vref vspike_down vres vdd
Xppolyf_u_resistor$3_20 vdd m1_132_n49# vspike_up ppolyf_u_resistor$3
Xppolyf_u_resistor$3_21 vdd m1_132_n49# vdd ppolyf_u_resistor$3
Xppolyf_u_resistor$3_10 vdd vref m1_600_n2985# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_11 vdd vref m1_n236_n2985# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_12 vdd vref m1_n236_n1981# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_13 vdd vref m1_600_n1981# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_14 vdd m1_56_n1479# m1_n236_n1981# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_15 vdd m1_308_n1479# m1_600_n1981# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_16 vdd m1_308_n1479# m1_n236_n977# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_17 vdd m1_56_n1479# m1_n236_n977# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_18 vdd m1_132_n551# vspike_up ppolyf_u_resistor$3
Xppolyf_u_resistor$3_19 vdd m1_132_n551# m1_n236_n977# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_0 vdd m1_308_n4993# vss ppolyf_u_resistor$3
Xppolyf_u_resistor$3_1 vdd m1_56_n4993# vss ppolyf_u_resistor$3
Xppolyf_u_resistor$3_2 vdd m1_308_n4993# m1_600_n4492# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_3 vdd m1_56_n4993# m1_n236_n4491# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_4 vdd vres m1_n236_n4491# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_5 vdd vres m1_600_n4492# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_6 vdd m1_132_n3563# vres ppolyf_u_resistor$3
Xppolyf_u_resistor$3_7 vdd m1_132_n3563# vspike_down ppolyf_u_resistor$3
Xppolyf_u_resistor$3_8 vdd vspike_down m1_600_n2985# ppolyf_u_resistor$3
Xppolyf_u_resistor$3_9 vdd vspike_down m1_n236_n2985# ppolyf_u_resistor$3
.ends

.subckt nfet$20 a_n256_n198# a_38_n60# a_n84_0# a_138_0#
X0 a_138_0# a_38_n60# a_n84_0# a_n256_n198# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$17 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$1$5 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$3$2 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt pfet$1$10 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt ota_1stage$2 vss vdd vp vn vout
Xnfet$17_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$17
Xnfet$17_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$17
Xnfet$1$5_0 vss vn vout m2_n516_n58# nfet$1$5
Xnfet$3$2_0 m2_n1824_n806# vss vdd vdd nfet$3$2
Xnfet$1$5_1 vss vp m2_n516_n58# m2_n346_983# nfet$1$5
Xpfet$1$10_0 pfet$1$10_1/w_n352_n286# vout vdd m2_n346_983# pfet$1$10
Xpfet$1$10_1 pfet$1$10_1/w_n352_n286# vdd m2_n346_983# m2_n346_983# pfet$1$10
.ends

.subckt ppolyf_u_resistor$2 a_n376_0# a_160_0# a_n132_0#
X0 a_n132_0# a_160_0# a_n376_0# ppolyf_u r_width=0.8u r_length=0.8u
.ends

.subckt pfet$18 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$24 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$3 vdd cntrl out in2 in1 m2_n850_n472# vss
Xpfet$18_2 m2_n850_n472# cntrl vdd vdd pfet$18
Xnfet$24_1 vss cntrl in2 out nfet$24
Xnfet$24_2 vss cntrl m2_n850_n472# vss nfet$24
Xpfet$18_0 out cntrl in1 vdd pfet$18
Xpfet$18_1 in2 m2_n850_n472# out vdd pfet$18
Xnfet$24_0 vss m2_n850_n472# out in1 nfet$24
.ends

.subckt nfet$22 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$17 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$23 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$21 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_1stage$3 vss vdd vp vn vout
Xnfet$22_0 vss vn vout m2_n516_n58# nfet$22
Xnfet$22_1 vss vp m2_n516_n58# m2_n346_983# nfet$22
Xpfet$17_0 pfet$17_1/w_n352_n286# vout vdd m2_n346_983# pfet$17
Xpfet$17_1 pfet$17_1/w_n352_n286# vdd m2_n346_983# m2_n346_983# pfet$17
Xnfet$23_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$23
Xnfet$23_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$23
Xnfet$21_0 m2_n1824_n806# vss vdd vdd nfet$21
>>>>>>> 32141c32e70fca95ef182d405dd80b0d5ace3811
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

<<<<<<< HEAD
.subckt pfet$26 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$42 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt switch out cntrl in vdd vss
Xpfet$26_0 m2_n331_n296# cntrl vdd vdd pfet$26
Xpfet$26_1 in m2_n331_n296# out vdd pfet$26
Xnfet$42_0 vss cntrl m2_n331_n296# vss nfet$42
Xnfet$42_1 vss cntrl in out nfet$42
.ends

.subckt nfet$47 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.3355p pd=2.32u as=0.3355p ps=2.32u w=0.55u l=0.28u
.ends

.subckt nfet$45 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$46 a_n256_n272# a_n84_0# a_198_0# a_38_n132#
X0 a_198_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.8u
.ends

.subckt nfet$44 a_n84_n2# a_n256_n272# a_30_n132# a_94_0#
X0 a_94_0# a_30_n132# a_n84_n2# a_n256_n272# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
.ends

.subckt nvdiv vss vdd vspike_up vspike_down vres vref
Xnfet$47_0 vss vdd vdd vref nfet$47
Xnfet$45_0 vss vspike_down vspike_down vres nfet$45
Xnfet$45_1 vss m2_367_1540# m2_367_1540# vspike_down nfet$45
Xnfet$46_0 vss vres vss vres nfet$46
Xnfet$44_0 vref vss vref vss nfet$44
Xnfet$44_1 vspike_up vss vspike_up m2_367_1540# nfet$44
Xnfet$44_2 vdd vss vdd vspike_up nfet$44
.ends

.subckt cap_mim$2 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt nfet$32 a_98_0# a_n256_n272# a_n84_0# a_32_n132#
X0 a_98_0# a_32_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
.ends

.subckt pfet$20 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$31 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt not$1 out in vdd vss
Xpfet$20_0 out in vdd vdd pfet$20
Xnfet$31_0 vss in out vss nfet$31
.ends

.subckt nfet$29 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$19 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$30 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$18 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nand$1 A B Z vdd vss
Xnfet$29_0 vss B nfet$30_0/a_94_0# vss nfet$29
Xpfet$19_0 B Z vdd vdd pfet$19
Xnfet$30_0 A Z nfet$30_0/a_94_0# vss nfet$30
Xpfet$18_0 A vdd vdd Z pfet$18
.ends

.subckt monostable vin vres vneg phi_1 phi_2 vss vdd
Xcap_mim$2_0 not$1_1/in nand$1_0/Z cap_mim$2
Xcap_mim$2_1 not$1_3/in nand$1_1/Z cap_mim$2
Xnfet$32_0 vss vss not$1_1/in vres nfet$32
Xnfet$32_1 vss vss not$1_3/in vres nfet$32
Xnot$1_0 phi_2 not$1_0/in vdd vss not$1
Xnot$1_1 not$1_0/in not$1_1/in vdd vss not$1
Xnot$1_2 phi_1 vneg vdd vss not$1
Xnot$1_3 vneg not$1_3/in vdd vss not$1
Xnand$1_0 not$1_0/in phi_1 nand$1_0/Z vdd vss nand$1
Xnand$1_1 vneg vin nand$1_1/Z vdd vss nand$1
.ends

.subckt pfet$23 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt pfet$24 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$39 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$40 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nor A B Z vdd vss
Xpfet$23_0 B vdd Z pfet$23_0/a_94_0# pfet$23
Xpfet$24_0 A pfet$23_0/a_94_0# vdd vdd pfet$24
Xnfet$39_0 vss A Z vss nfet$39
Xnfet$40_0 B vss Z vss nfet$40
.ends

.subckt nfet$43 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$27 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt conmutator out in1 in2 vdd cntrl vss
Xnfet$43_0 vss m2_n850_n472# out in1 nfet$43
Xnfet$43_2 vss cntrl m2_n850_n472# vss nfet$43
Xnfet$43_1 vss cntrl in2 out nfet$43
Xpfet$27_0 out cntrl in1 vdd pfet$27
Xpfet$27_1 in2 m2_n850_n472# out vdd pfet$27
Xpfet$27_2 m2_n850_n472# cntrl vdd vdd pfet$27
.ends

.subckt nfet$38 a_n256_n198# a_n84_0# a_94_0# a_30_1060#
X0 a_94_0# a_30_1060# a_n84_0# a_n256_n198# nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.28u
.ends

.subckt nfet$36 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$37 a_n84_n2# a_n256_n198# a_638_0# a_38_n60#
X0 a_638_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=3u
.ends

.subckt pfet$21 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$34 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$35 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$33 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_1stage$1 vdd vp vn vss vout
Xpfet$21_0 vdd vdd m3_n314_178# m3_n314_178# pfet$21
Xpfet$21_1 vdd vdd vout m3_n314_178# pfet$21
Xnfet$34_0 vss vn m3_n530_n14# vout nfet$34
Xnfet$34_1 vss vp m3_n530_n14# m3_n314_178# nfet$34
Xnfet$35_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$35
Xnfet$35_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$35
Xnfet$33_0 m3_n1200_n476# vss vdd vdd nfet$33
.ends

.subckt refractory vneg vspike_down vss vdd vrefrac
Xnfet$38_0 vss ota_1stage$1_0/vp vss ota_1stage$1_0/vp nfet$38
Xnfet$36_0 vss ota_1stage$1_0/vn vspike_down vspike_down nfet$36
Xnfet$36_1 vss vrefrac ota_1stage$1_0/vn ota_1stage$1_0/vn nfet$36
Xnfet$37_0 ota_1stage$1_0/vp vss vneg vneg nfet$37
Xota_1stage$1_0 vdd ota_1stage$1_0/vp ota_1stage$1_0/vn vss vrefrac ota_1stage$1
.ends

.subckt nfet$41 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$25 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt not$2 out in vdd vss
Xnfet$41_0 vss in out vss nfet$41
Xpfet$25_0 out in vdd vdd pfet$25
.ends

.subckt phaseUpulse phi_fire vin vres vspike reward vdd vref vss
Xswitch_0 switch_0/out phi_1 vspike vdd vss switch
Xswitch_1 vrefrac phi_2 vspike vdd vss switch
Xswitch_2 vref phi_int vspike vdd vss switch
Xnvdiv_0 vss vdd vspike_up vspike_down vres vref nvdiv
Xmonostable_0 vin vres vneg phi_1 phi_2 vss vdd monostable
Xnor_0 phi_1 phi_2 phi_int vdd vss nor
Xconmutator_0 switch_0/out vspike_up vdd vdd reward vss conmutator
Xrefractory_0 vneg vspike_down vss vdd vrefrac refractory
Xnot$2_0 phi_fire phi_int vdd vss not$2
.ends

.subckt LIF_comp vin vdd vss vout v_rew
Xota_1stage$2_0 vdd ota_1stage$2_0/vp v_th vss phaseUpulse_0/vin ota_1stage$2
Xnfet$50_0 vss v_th vin vmem nfet$50
Xota_2stage_0 vdd vspike vin vss vmem ota_2stage
Xswitch$1_0 vmem phi_fire vin vdd vss switch$1
Xconmutator$1_0 vmem vss vdd ota_1stage$2_0/vp phi_fire vss conmutator$1
Xcap_mim$3_0 conmutator$1_2/out vin cap_mim$3
Xconmutator$1_1 v_ref vmem vdd vout phi_fire vss conmutator$1
Xconmutator$1_2 vmem v_ref vdd conmutator$1_2/out phi_fire vss conmutator$1
XphaseUpulse_0 phi_fire phaseUpulse_0/vin v_th vspike v_rew vdd v_ref vss phaseUpulse
=======
.subckt nfet$15 a_n84_n2# a_238_0# a_n256_n272# a_38_n132#
X0 a_238_0# a_38_n132# a_n84_n2# a_n256_n272# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=1u
.ends

.subckt nfet$2$4 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$1$7 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$3$5 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$11 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nand$4 Z A B vdd vss
Xnfet$2$4_0 vss B nfet$3$5_0/a_94_0# vss nfet$2$4
Xpfet$1$7_0 B Z vdd vdd pfet$1$7
Xnfet$3$5_0 A Z nfet$3$5_0/a_94_0# vss nfet$3$5
Xpfet$11_0 A vdd vdd Z pfet$11
.ends

.subckt nfet$11 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$13 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt not$1 vss in out vdd
Xnfet$11_0 vss in out vss nfet$11
Xpfet$13_0 out in vdd vdd pfet$13
.ends

.subckt pfet$7 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$8 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt not vss vdd in
Xpfet$7_0 in in vdd vdd pfet$7
Xnfet$8_0 vss in in vss nfet$8
.ends

.subckt nfet$13 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$15 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt switch$1 vss out in cntrl vdd
Xnfet$13_0 vss cntrl m2_n331_n296# vss nfet$13
Xnfet$13_1 vss cntrl in out nfet$13
Xpfet$15_0 m2_n331_n296# cntrl vdd vdd pfet$15
Xpfet$15_1 in m2_n331_n296# out vdd pfet$15
.ends

.subckt pfet$1$8 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt pfet$2$7 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$10 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$1$3 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nor$2 B Z vdd m1_n7_n472# A vss
Xpfet$1$8_0 m1_n7_n472# vdd Z pfet$1$8_0/a_94_0# pfet$1$8
Xpfet$2$7_0 A pfet$1$8_0/a_94_0# vdd vdd pfet$2$7
Xnfet$10_0 vss A Z vss nfet$10
Xnfet$1$3_0 m1_n7_n472# vss Z vss nfet$1$3
.ends

.subckt nfet$16 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.915p pd=4.22u as=0.915p ps=4.22u w=1.5u l=0.28u
.ends

.subckt pfet$14 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$12 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$1 cntrl out in2 in1 vdd vss
Xpfet$14_0 out cntrl in1 vdd pfet$14
Xpfet$14_1 in2 m2_n850_n472# out vdd pfet$14
Xpfet$14_2 m2_n850_n472# cntrl vdd vdd pfet$14
Xnfet$12_0 vss m2_n850_n472# out in1 nfet$12
Xnfet$12_1 vss cntrl in2 out nfet$12
Xnfet$12_2 vss cntrl m2_n850_n472# vss nfet$12
.ends

.subckt nfet$8$1 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt phaseUpulse reward phi_int vin vspike m4_n522_1747# m2_2886_n700# nand$4_0/Z
+ a_1700_n1729# not$1_0/out m4_1944_1747# vspike_up m2_1332_n780# switch$1_1/in not_3/vdd
+ m1_2078_n924# switch$1_2/in not_3/vss phi_2 nand$4_1/Z vneg
Xnfet$15_0 m2_554_n1578# vneg not_3/vss m2_554_n1578# nfet$15
Xnand$4_0 nand$4_0/Z vin vneg not_3/vdd not_3/vss nand$4
Xnand$4_1 nand$4_1/Z vneg phi_2 not_3/vdd not_3/vss nand$4
Xnot$1_0 not_3/vss phi_int not$1_0/out not_3/vdd not$1
Xnot_0 not_3/vss not_3/vdd vneg not
Xswitch$1_0 not_3/vss vspike switch$1_0/in vneg not_3/vdd switch$1
Xnot_1 not_3/vss not_3/vdd vneg not
Xnor$2_0 nor$2_0/B phi_int not_3/vdd vneg phi_2 not_3/vss nor$2
Xnot_2 not_3/vss not_3/vdd phi_2 not
Xswitch$1_1 not_3/vss vspike switch$1_1/in phi_2 not_3/vdd switch$1
Xnfet$16_0 not_3/vss not_3/vss not_3/vss m2_554_n1578# nfet$16
Xswitch$1_2 not_3/vss vspike switch$1_2/in phi_int not_3/vdd switch$1
Xnot_3 not_3/vss not_3/vdd phi_2 not
Xconmutator$1_0 reward vspike not_3/vdd vspike_up not_3/vdd not_3/vss conmutator$1
Xnfet$8$1_0 not_3/vss m1_2078_n924# m1_2078_n924# m2_1332_n780# nfet$8$1
Xnfet$8$1_2 not_3/vss m4_n522_1747# m2_n103_1601# not_3/vss nfet$8$1
Xnfet$8$1_1 not_3/vss m1_2078_n924# m2_2886_n700# m2_2886_n700# nfet$8$1
Xnfet$8$1_3 not_3/vss m4_1944_1747# m2_n103_1601# not_3/vss nfet$8$1
.ends

.subckt nfet$29 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt nfet$27 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$19 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt cap_mim$5 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt pfet$20 a_28_n136# a_n92_0# a_94_0# w_n352_n362#
X0 a_94_0# a_28_n136# a_n92_0# w_n352_n362# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
.ends

.subckt nfet$28 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$26 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_2stages$1 vss vdd vn vp pfet$20_0/w_n352_n362# vout
Xnfet$29_0 vss m2_n516_n58# vss vout nfet$29
Xnfet$27_0 vss vp m2_196_146# m2_n516_n58# nfet$27
Xnfet$27_1 vss vn m2_n516_n58# m2_n346_983# nfet$27
Xpfet$19_0 pfet$20_0/w_n352_n362# m2_196_146# vdd m2_n346_983# pfet$19
Xpfet$19_1 pfet$20_0/w_n352_n362# vdd m2_n346_983# m2_n346_983# pfet$19
Xcap_mim$5_0 vout m2_196_146# cap_mim$5
Xpfet$20_0 m2_196_146# vdd vout pfet$20_0/w_n352_n362# pfet$20
Xnfet$28_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$28
Xnfet$28_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$28
Xnfet$26_0 m2_n1824_n806# vss vdd vdd nfet$26
.ends

.subckt LIF_comp vout
Xcap_mim$4_0 phaseUpulse_0/phi_2 phaseUpulse_0/nand$4_1/Z cap_mim$4
Xvdiv$1_0 vdiv$1_0/vss vdiv$1_0/vspike_up vdiv$1_0/vref vdiv$1_0/vspike_down vdiv$1_0/vres
+ vdiv$1_0/vss vdiv$1
Xcap_mim$4_1 phaseUpulse_0/vneg phaseUpulse_0/nand$4_0/Z cap_mim$4
Xnfet$20_0 vdiv$1_0/vss ota_1stage$2_0/vn ota_2stages$1_0/vn conmutator$3_0/in1 nfet$20
Xota_1stage$2_0 vdiv$1_0/vss ota_1stage$2_0/vdd ota_1stage$2_0/vp ota_1stage$2_0/vn
+ phaseUpulse_0/vin ota_1stage$2
Xppolyf_u_resistor$2_0 vdiv$1_0/vss ota_1stage$2_0/vn vdiv$1_0/vss ppolyf_u_resistor$2
Xppolyf_u_resistor$2_1 vdiv$1_0/vss ota_1stage$2_0/vn m1_2167_4433# ppolyf_u_resistor$2
Xppolyf_u_resistor$2_2 vdiv$1_0/vss vdiv$1_0/vss m1_2167_4433# ppolyf_u_resistor$2
Xppolyf_u_resistor$2_3 vdiv$1_0/vss vdiv$1_0/vss ppolyf_u_resistor$2_3/a_n132_0# ppolyf_u_resistor$2
Xppolyf_u_resistor$2_4 vdiv$1_0/vss ota_1stage$2_0/vn vdiv$1_0/vss ppolyf_u_resistor$2
Xconmutator$3_0 vdiv$1_0/vss conmutator$3_0/cntrl ota_1stage$2_0/vp vdiv$1_0/vss conmutator$3_0/in1
+ conmutator$3_0/m2_n850_n472# vdiv$1_0/vss conmutator$3
Xconmutator$3_2 conmutator$3_2/vdd vdiv$1_0/vref conmutator$3_2/out conmutator$3_2/in2
+ conmutator$3_2/in1 conmutator$3_2/m2_n850_n472# vdiv$1_0/vss conmutator$3
Xconmutator$3_1 vdiv$1_0/vss conmutator$3_1/cntrl conmutator$3_1/out conmutator$3_1/in2
+ conmutator$3_1/in1 vout vdiv$1_0/vss conmutator$3
Xota_1stage$3_0 vdiv$1_0/vss vdiv$1_0/vss ota_1stage$3_0/vp ota_1stage$3_0/vn ota_1stage$3_0/vout
+ ota_1stage$3
Xcap_mim$3_0 vdiv$1_0/vref ota_2stages$1_0/vn cap_mim$3
XphaseUpulse_0 phaseUpulse_0/reward phaseUpulse_0/phi_int phaseUpulse_0/vin phaseUpulse_0/vspike
+ phaseUpulse_0/vneg vdiv$1_0/vspike_down phaseUpulse_0/nand$4_0/Z vdiv$1_0/vss conmutator$3_0/cntrl
+ phaseUpulse_0/phi_2 vdiv$1_0/vspike_up ota_1stage$3_0/vout vdiv$1_0/vref vdiv$1_0/vss
+ ota_1stage$3_0/vn ota_1stage$3_0/vout vdiv$1_0/vss phaseUpulse_0/phi_2 phaseUpulse_0/nand$4_1/Z
+ phaseUpulse_0/vneg phaseUpulse
Xota_2stages$1_0 vdiv$1_0/vss vdiv$1_0/vss ota_2stages$1_0/vn ota_2stages$1_0/vp w_954_1524#
+ conmutator$3_0/in1 ota_2stages$1
>>>>>>> 32141c32e70fca95ef182d405dd80b0d5ace3811
.ends

