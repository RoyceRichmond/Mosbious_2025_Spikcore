* NGSPICE file created from AH_neuron.ext - technology: gf180mcuD

.subckt pfet a_38_n60# a_n92_0# a_318_0# w_n230_n138#
X0 a_318_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=1.4u
.ends

.subckt nfet$7 a_n84_n2# a_374_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_374_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=1.68u
.ends

.subckt nfet a_150_0# dw_n710_n726# a_n84_0# a_38_n132# w_n710_n726#
X0 a_150_0# a_38_n132# a_n84_0# w_n710_n726# nfet_03v3 ad=0.2684p pd=2.1u as=0.2684p ps=2.1u w=0.44u l=0.56u
.ends

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=6u c_length=5u
.ends

.subckt nfet$6 a_1158_0# a_n84_n2# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_1158_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=5.6u
.ends

.subckt pfet$1 a_150_0# a_38_n60# a_n92_0# w_n230_n138#
X0 a_150_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.286p pd=2.18u as=0.286p ps=2.18u w=0.44u l=0.56u
.ends

.subckt nfet$4 a_n84_n2# a_194_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_194_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.78u
.ends

.subckt AH_neuron vdd Current_in v_bias vss vout
Xpfet_0 m2_381_1901# vout vdd vdd pfet
Xnfet$7_0 m1_335_n170# vss nfet_0/dw_n710_n726# vout vss nfet$7
Xnfet_0 vss nfet_0/dw_n710_n726# m2_381_1901# Current_in vss nfet
Xcap_mim$1_0 Current_in vout cap_mim$1
Xnfet$6_0 m1_335_n170# Current_in nfet_0/dw_n710_n726# v_bias vss nfet$6
Xpfet$1_0 vdd Current_in m2_381_1901# vdd pfet$1
Xnfet$4_0 vout vss nfet_0/dw_n710_n726# m2_381_1901# vss nfet$4
.ends

