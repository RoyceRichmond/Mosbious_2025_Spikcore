magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
rect 0 0 1 1
<< l46d0 >>
rect 0 0 1 1
<< l41d0 >>
<< l81d0 >>
rect 0 0 1 1
<< l117d5 >>
rect 0 0 1 1
<< l117d10 >>
<< l75d0 >>
rect 0 0 1 1
<< labels >>
rlabel l81d10 0.25 0.25 0.25 0.25 0 
rlabel l46d10 0.25 -0.03 0.25 -0.03 0 
<< end >>
