magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
rect 0 0 4 4
<< l34d0 >>
<< l36d0 >>
<< l42d0 >>
rect 1 1 2 2
<< l81d0 >>
rect 3 1 4 4
<< labels >>
rlabel l34d10 3.3725 0.648 3.3725 0.648 0 vss
rlabel l34d10 3.112 0.846 3.112 0.846 0 phi_fire
rlabel l34d10 0.087 0.928 0.087 0.928 0 vin
rlabel l42d10 1.8865 1.8475 1.8865 1.8475 0 vrefrac
rlabel l42d10 2.798 1.1645 2.798 1.1645 0 phi_int
rlabel l42d10 2.2565 1.1675 2.2565 1.1675 0 phi_2
rlabel l42d10 1.4995 1.1665 1.4995 1.1665 0 phi_1
rlabel l42d10 2.5495 1.8515 2.5495 1.8515 0 vref
rlabel l42d10 0.9225 1.206 0.9225 1.206 0 vneg
rlabel l81d10 3.5065 3.885 3.5065 3.885 0 vss
rlabel l81d10 3.626 3.8765 3.626 3.8765 0 vdd
rlabel l36d10 1.738 1.346 1.738 1.346 0 vspike
rlabel l36d10 0.746 1.532 0.746 1.532 0 reward
rlabel l36d10 0.4275 3.2795 0.4275 3.2795 0 vspike_up
rlabel l36d10 0.8765 3.3765 0.8765 3.3765 0 vspike_down
rlabel l36d10 1.154 3.19 1.154 3.19 0 vres
rlabel l36d10 2.9355 0.8585 2.9355 0.8585 0 phi_int
use monostable monostable_1
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 3 2
use refractory refractory_1
timestamp 1757365861
transform -1 0 2 0 1 2
box -1 -1 1 1
use vdiv vdiv_1
timestamp 1757365861
transform -1 0 3 0 -1 4
box 0 0 2 1
use nor nor_1
timestamp 1757365861
transform -1 0 3 0 1 1
box 0 0 0 0
use notx241 notx241_1
timestamp 1757365861
transform -1 0 3 0 1 1
box 0 0 0 0
use via_devx2424x241 via_devx2424x241_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2424x241 via_devx2424x241_2
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_2
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2426x241 via_devx2426x241_1
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2426x241 via_devx2426x241_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2426x241 via_devx2426x241_3
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2426x241 via_devx2426x241_4
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use switch switch_1
timestamp 1757365861
transform 1 0 3 0 -1 1
box 0 0 0 0
use conmutator conmutator_1
timestamp 1757365861
transform 1 0 1 0 -1 1
box -1 0 0 0
use via_devx2425x241 via_devx2425x241_3
timestamp 1757365861
transform 1 0 3 0 1 2
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_4
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use switch switch_2
timestamp 1757365861
transform 1 0 2 0 -1 1
box 0 0 0 0
use via_devx2424x241 via_devx2424x241_3
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_5
timestamp 1757365861
transform 1 0 2 0 1 2
box 0 0 0 0
use switch switch_3
timestamp 1757365861
transform 1 0 1 0 -1 1
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_6
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2425x241 via_devx2425x241_7
timestamp 1757365861
transform 1 0 1 0 1 2
box 0 0 0 0
use via_devx2432 via_devx2432_1
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2432 via_devx2432_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2432 via_devx2432_3
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2432 via_devx2432_4
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2433 via_devx2433_1
timestamp 1757365861
transform 1 0 2 0 1 2
box 0 0 0 0
use via_devx2433 via_devx2433_2
timestamp 1757365861
transform 1 0 1 0 1 2
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2434 via_devx2434_1
timestamp 1757365861
transform 1 0 3 0 1 2
box 0 0 0 0
use via_devx2433 via_devx2433_3
timestamp 1757365861
transform 1 0 3 0 1 3
box 0 0 0 0
use via_devx2432 via_devx2432_5
timestamp 1757365861
transform 1 0 2 0 1 3
box 0 0 0 0
use via_devx2433 via_devx2433_4
timestamp 1757365861
transform 1 0 1 0 1 2
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_2
timestamp 1757365861
transform 1 0 1 0 1 3
box 0 0 0 0
use via_devx2433 via_devx2433_5
timestamp 1757365861
transform 1 0 0 0 1 2
box 0 0 0 0
use via_devx2432 via_devx2432_6
timestamp 1757365861
transform 1 0 3 0 1 3
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_3
timestamp 1757365861
transform 1 0 0 0 1 3
box 0 0 0 0
use via_devx2432 via_devx2432_7
timestamp 1757365861
transform 1 0 2 0 1 3
box 0 0 0 0
use via_devx2433 via_devx2433_6
timestamp 1757365861
transform 1 0 2 0 1 0
box 0 0 0 0
use via_devx2432 via_devx2432_8
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_4
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_5
timestamp 1757365861
transform 1 0 1 0 1 3
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_6
timestamp 1757365861
transform 1 0 2 0 1 0
box 0 0 0 0
use via_devx2432x241 via_devx2432x241_7
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use via_devx2434x241 via_devx2434x241_1
timestamp 1757365861
transform 1 0 3 0 1 4
box 0 0 0 0
use via_devx2434x241 via_devx2434x241_2
timestamp 1757365861
transform 1 0 3 0 1 2
box 0 0 0 0
use via_devx2434x241 via_devx2434x241_3
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2434x241 via_devx2434x241_4
timestamp 1757365861
transform 1 0 4 0 1 3
box 0 0 0 0
use via_devx2434x241 via_devx2434x241_5
timestamp 1757365861
transform 1 0 4 0 1 1
box 0 0 0 0
<< end >>
