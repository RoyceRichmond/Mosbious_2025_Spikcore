* Extracted by KLayout with GF180 LVS runset on : 09/08/2025 07:51

.SUBCKT DFF_2phase_1 D PHI_1 PHI_2 out_m Q gf180mcu_gnd
X$1 \$7 out_m PHI_1 D \$6 \$6 gf180mcu_gnd gf180mcu_fd_sc_mcu9t5v0__latq_1
X$4 \$7 Q PHI_2 out_m \$6 \$6 gf180mcu_gnd gf180mcu_fd_sc_mcu9t5v0__latq_1
.ENDS DFF_2phase_1

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__latq_1 VSS Q E D VDD \$21 gf180mcu_gnd
M$1 VDD \$4 Q \$21 pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$2 \$17 D VDD \$21 pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$3 \$4 \$2 \$17 \$21 pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U PD=1.52U
M$4 \$4 \$3 \$18 \$21 pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U PD=1.52U
M$5 VDD \$5 \$18 \$21 pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$6 \$5 \$4 VDD \$21 pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$7 VDD E \$2 \$21 pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$8 \$3 \$2 VDD \$21 pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U PD=2.88U
M$9 VSS \$4 Q gf180mcu_gnd nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$10 \$10 D VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$11 \$4 \$3 \$10 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$12 \$9 \$2 \$4 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$13 VSS \$5 \$9 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$14 \$5 \$4 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$15 VSS E \$2 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$16 \$3 \$2 VSS gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
.ENDS gf180mcu_fd_sc_mcu9t5v0__latq_1
