** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/pex/LIF_ring/LIF_ring.sch
**.subckt LIF_ring vdd vlk vout vss
V1 net2 GND 1.8
Vdd_c net3 vdd 0
.save i(vdd_c)
R1 net3 net2 10 m=1
V2 net1 GND 0.2
x1 vdd net1 spk GND LIF_ring
**** begin user architecture code


.option method=gear seed=12
.tran 0.01n 5u
.include /foss/designs/Mosbious_2025_Spikcore/designs/pex/LIF_ring/LIF_ring_pex.spice
.save allcurrents
.options save currents
.control
	reset
	save all
        run
        write LIF_ring.raw
.endc



.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
