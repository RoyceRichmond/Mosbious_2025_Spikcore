magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
rect 0 0 2 1
<< l34d0 >>
<< labels >>
rlabel l34d10 0.5435 0.534 0.5435 0.534 0 vdd
rlabel l34d10 0.595 -0.276 0.595 -0.276 0 vss
rlabel l34d10 0.1695 0.001 0.1695 0.001 0 vspike_up
rlabel l34d10 0.6295 0.002 0.6295 0.002 0 vref
rlabel l34d10 1.1075 0.106 1.1075 0.106 0 vspike_down
rlabel l34d10 1.5935 0.261 1.5935 0.261 0 vres
use ppolyf_u_resistor ppolyf_u_resistor_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx241 ppolyf_u_resistorx241_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx242 ppolyf_u_resistorx242_1
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx242 ppolyf_u_resistorx242_2
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx243 ppolyf_u_resistorx243_1
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx241 ppolyf_u_resistorx241_2
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx244 ppolyf_u_resistorx244_1
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use ppolyf_u_resistorx242 ppolyf_u_resistorx242_3
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
<< end >>
