* NGSPICE file created from refractory.ext - technology: gf180mcuD

.subckt pfet w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$1 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt nfet$2 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt ota_1stage vdd vp vn vss vout
Xpfet_0 vdd vdd m3_n314_178# m3_n314_178# pfet
Xpfet_1 vdd vdd vout m3_n314_178# pfet
Xnfet$1_0 vss vn m3_n530_n14# vout nfet$1
Xnfet$1_1 vss vp m3_n530_n14# m3_n314_178# nfet$1
Xnfet_0 m3_n1200_n476# vss vdd vdd nfet
Xnfet$2_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$2
Xnfet$2_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$2
.ends

.subckt nfet$3 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$6 a_n84_n2# a_n256_n198# a_638_0# a_38_n60#
X0 a_638_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=3u
.ends

.subckt nfet$4 a_n256_n198# a_n84_0# a_94_0# a_30_1060#
X0 a_94_0# a_30_1060# a_n84_0# a_n256_n198# nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.28u
.ends

.subckt refractory vneg vspike_down vss vdd vrefrac
Xota_1stage_0 vdd ota_1stage_0/vp ota_1stage_0/vn vss vrefrac ota_1stage
Xnfet$3_0 vss ota_1stage_0/vn vspike_down vspike_down nfet$3
Xnfet$3_1 vss vrefrac ota_1stage_0/vn ota_1stage_0/vn nfet$3
Xnfet$6_0 ota_1stage_0/vp vss vneg vneg nfet$6
Xnfet$4_0 vss ota_1stage_0/vp vss ota_1stage_0/vp nfet$4
.ends

