** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/klayout/layout_top/top.sch
.subckt top PIN[15] PIN[16] PIN[17] PIN[18] PIN[19] PIN[20] PIN[21] PIN[22] VDD VSS PIN[1] PIN[2] V_EX V_INH PIN[3] PIN[4]
+ PIN[5] PIN[6] PIN[7] PIN[8] EN DATA CLK PIN[23] PIN[24] PIN[9] PIN[10] PIN[11] PIN[12] PIN[13] PIN[14] VAH_bias
*.PININFO PIN[15]:B PIN[16]:B PIN[17]:B PIN[18]:B PIN[19]:B PIN[20]:B PIN[21]:B PIN[22]:B VDD:B VSS:B PIN[1]:B PIN[2]:B V_EX:B
*+ V_INH:B PIN[3]:B PIN[4]:B PIN[5]:B PIN[6]:B PIN[7]:B PIN[8]:B EN:B DATA:B CLK:B PIN[23]:B PIN[24]:B PIN[9]:B PIN[10]:B PIN[11]:B
*+ PIN[12]:B PIN[13]:B PIN[14]:B VAH_bias:B
x5 VDD VSS PIN[1] VSS PIN[2] LIF_comp
x6 VDD PIN[3] V_EX net1 PIN[4] V_INH VSS synapse
x2 VDD PIN[5] V_EX net2 PIN[6] V_INH VSS synapse
x3 VDD PIN[7] V_EX net3 PIN[8] V_INH VSS synapse
x7 VDD PIN[9] V_EX net4 PIN[10] V_INH VSS synapse
x8 VDD PIN[11] V_EX net5 PIN[12] V_INH VSS synapse
x9 VDD PIN[13] V_EX net6 PIN[14] V_INH VSS synapse
x10 VDD PIN[15] PIN[16] VSS VAH_bias AH_neuron
x11 VDD PIN[17] PIN[18] VSS VAH_bias AH_neuron
x12 VDD PIN[19] PIN[20] VSS VAH_bias AH_neuron
x13 VDD PIN[21] PIN[22] VSS VAH_bias AH_neuron
x14 VDD PIN[23] PIN[24] VSS VAH_bias AH_neuron
x1 clk_schmitt CLK VDD VSS schmitt_trigger
x4 data_schmitt DATA VDD VSS schmitt_trigger
x15 net7 net8 net8 net8 net8 net8 net8 net8 net8 net8 net8 PIN[1] PIN[2] PIN[3] PIN[4] PIN[5] PIN[6] PIN[7] PIN[8] PIN[9] PIN[10]
+ PIN[11] PIN[12] PIN[13] PIN[14] PIN[15] PIN[16] PIN[17] PIN[18] PIN[19] PIN[20] PIN[21] PIN[22] PIN[23] PIN[24] data_schmitt VDD EN
+ VSS clk_schmitt swmatrix_24_by_10
* noconn #net7
* noconn #net8
.ends

* expanding   symbol:  designs/libs/core_LIF_comp/LIF_comp.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/LIF_comp.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/LIF_comp.sch
.subckt LIF_comp vdd vss vin v_rew vout
*.PININFO vin:B v_rew:B vdd:B vss:B vout:B
x8 phi_fire vdd v_ref net1 vmem vss conmutator
x9 vdd v_ocomp v_icomp v_th vss ota_1stage
x10 vdd vin vmem vspike vss ota_2stage
x11 vdd vin vmem phi_fire vss switch
x12 phi_fire vdd vmem vout v_ref vss conmutator
x13 phi_fire vdd vss v_icomp vmem vss conmutator
x14 vss vdd v_ocomp vspike phi_fire v_ref v_rew v_th phaseUpulse
XC1 vin net1 cap_mim_2f0fF c_width=9e-6 c_length=9e-6 m=1
XM2 vmem v_th vin vss nfet_03v3 L=0.5u W=0.5u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_synapse/synapse.sym # of pins=7
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_synapse/synapse.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_synapse/synapse.sch
.subckt synapse vdd v_in ve v_ctrl v_out vi vss
*.PININFO v_out:B v_ctrl:B ve:B vi:B v_in:B vdd:B vss:B
XM5 net2 net2 vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM1 net1 v_in vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM3 net1 v_in vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM4 net2 v_in net3 vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM6 net3 ve vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM7 net5 vi vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM8 net4 net1 net5 vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM9 net4 net4 vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM2 net7 net2 vdd vdd pfet_03v3 L=0.28u W=2.8u nf=1 m=1
XM10 v_out v_ctrl net7 vdd pfet_03v3 L=0.28u W=2.8u nf=1 m=1
XM11 v_out v_ctrl net6 vss nfet_03v3 L=0.28u W=2u nf=1 m=1
XM12 net6 net4 vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_AH_neuron/AH_neuron.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_AH_neuron/AH_neuron.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_AH_neuron/AH_neuron.sch
.subckt AH_neuron vdd Current_in vout vss v_bias
*.PININFO vdd:B vss:B Current_in:B vout:B v_bias:B
XM5 vout net1 vdd vdd pfet_03v3 L=1.4u W=0.84u nf=1 m=1
XM1 net1 Current_in vdd vdd pfet_03v3 L=0.56u W=0.44u nf=1 m=1
XM2 vout net1 vss vss nfet_03v3 L=0.78u W=0.42u nf=1 m=1
XM3 net1 Current_in vss vss nfet_03v3 L=0.56u W=0.44u nf=1 m=1
XM4 net2 vout vss vss nfet_03v3 L=1.68u W=0.42u nf=1 m=1
XC3 vout Current_in cap_mim_2f0fF c_width=6e-6 c_length=5e-6 m=1
XM6 Current_in v_bias net2 vss nfet_03v3 L=5.6u W=0.42u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_schmitt_trigger/schmitt_trigger.sym # of pins=4
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_schmitt_trigger/schmitt_trigger.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_schmitt_trigger/schmitt_trigger.sch
.subckt schmitt_trigger out in vdd vss
*.PININFO in:I out:O vdd:B vss:B
XM2 outx in vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XM1 outz in vss vss nfet_03v3 L=0.28u W=2.1u nf=1 m=1
XM4 outy in outz vss nfet_03v3 L=0.28u W=2u nf=1 m=1
XM3 outx in outy vss nfet_03v3 L=0.28u W=2.5u nf=1 m=1
XM5 vdd outy outz vss nfet_03v3 L=0.28u W=1.1u nf=1 m=1
XM6 vdd outx outy vss nfet_03v3 L=0.3u W=1u nf=1 m=1
XM8 out outx vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM7 out outx vdd vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
XM10 outy vss vdd vdd pfet_03v3 L=0.8u W=1.6u nf=1 m=1
XM11 outx vss vdd vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
XM12 outy vdd vss vss nfet_03v3 L=2u W=0.42u nf=1 m=1
XM13 outx vdd vss vss nfet_03v3 L=0.6u W=1u nf=1 m=1
XM19 outz outz vdd vdd pfet_03v3 L=0.28u W=0.8u nf=1 m=1
XM15 outx out vdd vdd pfet_03v3 L=1u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_24_10/swmatrix_24_by_10.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_24_10/swmatrix_24_by_10.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_24_10/swmatrix_24_by_10.sch
.subckt swmatrix_24_by_10 D_out BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1] PIN[2] PIN[3] PIN[4]
+ PIN[5] PIN[6] PIN[7] PIN[8] PIN[9] PIN[10] PIN[11] PIN[12] PIN[13] PIN[14] PIN[15] PIN[16] PIN[17] PIN[18] PIN[19] PIN[20] PIN[21]
+ PIN[22] PIN[23] PIN[24] D_in VDD enable VSS clk
*.PININFO PIN[1:24]:B BUS[1:10]:B D_in:I D_out:O VDD:B VSS:B enable:I clk:B
xswmatrix_row[1] D_out_row[1] Data_in phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ VDD PIN[1] VSS swmatrix_row_10
xswmatrix_row[2] D_out_row[2] D_out_row[1] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[2] VSS swmatrix_row_10
xswmatrix_row[3] D_out_row[3] D_out_row[2] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[3] VSS swmatrix_row_10
xswmatrix_row[4] D_out_row[4] D_out_row[3] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[4] VSS swmatrix_row_10
xswmatrix_row[5] D_out_row[5] D_out_row[4] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[5] VSS swmatrix_row_10
xswmatrix_row[6] D_out_row[6] D_out_row[5] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[6] VSS swmatrix_row_10
xswmatrix_row[7] D_out_row[7] D_out_row[6] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[7] VSS swmatrix_row_10
xswmatrix_row[8] D_out_row[8] D_out_row[7] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[8] VSS swmatrix_row_10
xswmatrix_row[9] D_out_row[9] D_out_row[8] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[9] VSS swmatrix_row_10
xswmatrix_row[10] D_out_row[10] D_out_row[9] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[10] VSS swmatrix_row_10
xswmatrix_row[11] D_out_row[11] D_out_row[10] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[11] VSS swmatrix_row_10
xswmatrix_row[12] D_out_row[12] D_out_row[11] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[12] VSS swmatrix_row_10
xswmatrix_row[13] D_out_row[13] D_out_row[12] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[13] VSS swmatrix_row_10
xswmatrix_row[14] D_out_row[14] D_out_row[13] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[14] VSS swmatrix_row_10
xswmatrix_row[15] D_out_row[15] D_out_row[14] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[15] VSS swmatrix_row_10
xswmatrix_row[16] D_out_row[16] D_out_row[15] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[16] VSS swmatrix_row_10
xswmatrix_row[17] D_out_row[17] D_out_row[16] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[17] VSS swmatrix_row_10
xswmatrix_row[18] D_out_row[18] D_out_row[17] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[18] VSS swmatrix_row_10
xswmatrix_row[19] D_out_row[19] D_out_row[18] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[19] VSS swmatrix_row_10
xswmatrix_row[20] D_out_row[20] D_out_row[19] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[20] VSS swmatrix_row_10
xswmatrix_row[21] D_out_row[21] D_out_row[20] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[21] VSS swmatrix_row_10
xswmatrix_row[22] D_out_row[22] D_out_row[21] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[22] VSS swmatrix_row_10
xswmatrix_row[23] D_out_row[23] D_out_row[22] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9]
+ BUS[10] VDD PIN[23] VSS swmatrix_row_10
xswmatrix_row[24] D_out D_out_row[23] phi_1 phi_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ VDD PIN[24] VSS swmatrix_row_10
x1 phi_2 clock phi_1 VDD VSS NO_ClkGen
x4 VDD VSS clk clock enable D_in Data_in En_clk_din
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_conmutator/conmutator.sym # of pins=6
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_conmutator/conmutator.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_conmutator/conmutator.sch
.subckt conmutator cntrl vdd in2 out in1 vss
*.PININFO vdd:B vss:B in2:B out:B in1:B cntrl:B
x1 vdd cntrl net1 vss not
XM3 out net1 in2 vdd pfet_03v3 L=0.35u W=1u nf=1 m=1
XM4 out cntrl in2 vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM1 out cntrl in1 vdd pfet_03v3 L=0.35u W=1u nf=1 m=1
XM2 out net1 in1 vss nfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_ota_1stage/ota_1stage.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_ota_1stage/ota_1stage.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_ota_1stage/ota_1stage.sch
.subckt ota_1stage vdd vout vp vn vss
*.PININFO vdd:B vss:B vp:B vn:B vout:B
XM1 net1 net1 vdd vdd pfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM2 net1 vp net2 vss nfet_03v3 L=0.28u W=3.08u nf=1 m=1
XM4 vout net1 vdd vdd pfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM3 vout vn net2 vss nfet_03v3 L=0.28u W=3.08u nf=1 m=1
XM5 net2 net3 vss vss nfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM6 net3 net3 vss vss nfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM7 vdd vdd net3 vss nfet_03v3 L=8.54u W=0.36u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_ota_2stage/ota_2stage.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_ota_2stage/ota_2stage.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_ota_2stage/ota_2stage.sch
.subckt ota_2stage vdd vn vout vp vss
*.PININFO vdd:B vss:B vn:B vp:B vout:B
XM3 net1 net1 vdd vdd pfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM1 net1 vn net3 vss nfet_03v3 L=0.28u W=3.08u nf=1 m=1
XM4 net2 net1 vdd vdd pfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM2 net2 vp net3 vss nfet_03v3 L=0.28u W=3.08u nf=1 m=1
XM5 net3 net4 vss vss nfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM8 net4 net4 vss vss nfet_03v3 L=0.28u W=0.84u nf=1 m=1
XM9 vdd vdd net4 vss nfet_03v3 L=8.54u W=0.36u nf=1 m=1
XM6 vout net2 vdd vdd pfet_03v3 L=0.28u W=0.28u nf=1 m=6
XM7 vout net4 vss vss nfet_03v3 L=0.28u W=0.56u nf=1 m=1
XC1 net2 vout cap_mim_2f0fF c_width=9e-6 c_length=9e-6 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_switch/switch.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_switch/switch.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_switch/switch.sch
.subckt switch vdd in out cntrl vss
*.PININFO vdd:B vss:B in:B out:B cntrl:B
x1 vdd cntrl net1 vss not
XM3 out net1 in vdd pfet_03v3 L=0.35u W=1u nf=1 m=1
XM4 out cntrl in vss nfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_phaseUpulse/phaseUpulse.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_phaseUpulse/phaseUpulse.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_phaseUpulse/phaseUpulse.sch
.subckt phaseUpulse vss vdd vin vspike phi_fire vref reward vres
*.PININFO vin:I vdd:B vss:B vspike:O phi_fire:O vref:O reward:I vres:O
x19 vdd phi_int phi_fire vss not
x21 vdd vss phi_1 phi_2 phi_int nor
x7 vdd vspike net1 phi_1 vss switch
x10 vdd vspike vref phi_int vss switch
x18 vdd vspike vrefrac phi_2 vss switch
x20 reward vdd vdd net1 vspike_up vss conmutator
x6 vss vdd vin vres phi_1 phi_2 vneg monostable
x1 vss vdd vspike_down vneg vrefrac refractory
x2 vss vdd vref vspike_up vspike_down vres nvdiv
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_row_10/swmatrix_row_10.sym # of pins=9
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_row_10/swmatrix_row_10.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_row_10/swmatrix_row_10.sch
.subckt swmatrix_row_10 D_out D_in PHI_1 PHI_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] VDD
+ pin VSS
*.PININFO pin:B PHI_2:I PHI_1:I BUS[1:10]:B D_in:I D_out:O VDD:B VSS:B enable:I
xSR D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] D_out gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8] gc[9] gc[10] PHI_1
+ PHI_2 enable VDD VSS ShiftReg_row_10_2
xTgates[1] gc[1] BUS[1] pin VSS VDD swmatrix_Tgate
xTgates[2] gc[2] BUS[2] pin VSS VDD swmatrix_Tgate
xTgates[3] gc[3] BUS[3] pin VSS VDD swmatrix_Tgate
xTgates[4] gc[4] BUS[4] pin VSS VDD swmatrix_Tgate
xTgates[5] gc[5] BUS[5] pin VSS VDD swmatrix_Tgate
xTgates[6] gc[6] BUS[6] pin VSS VDD swmatrix_Tgate
xTgates[7] gc[7] BUS[7] pin VSS VDD swmatrix_Tgate
xTgates[8] gc[8] BUS[8] pin VSS VDD swmatrix_Tgate
xTgates[9] gc[9] BUS[9] pin VSS VDD swmatrix_Tgate
xTgates[10] gc[10] BUS[10] pin VSS VDD swmatrix_Tgate
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/NO_ClkGen/NO_ClkGen.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/NO_ClkGen/NO_ClkGen.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/NO_ClkGen/NO_ClkGen.sch
.subckt NO_ClkGen PHI_2 CLK PHI_1 VDD VSS
*.PININFO CLK:I PHI_2:O PHI_1:O VDD:B VSS:B
x1 OUT_bot_d CLKB OUT_top VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
x2 OUT_top_d CLKbuf OUT_bot VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
x3 OUT_top PHI_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x4 PHI_2 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x5 net3 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x6 OUT_bot PHI_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x7 PHI_1 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x8 net4 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x9 CLKB CLKbuf VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x10 CLK CLKB VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x11 net5 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x12 net6 net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x13 net2 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x15 net1 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x17 net7 net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x18 net8 net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x14 net9 net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x16 net12 net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x19 net10 OUT_top_d VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x20 net11 OUT_bot_d VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
* noconn VDD
* noconn VSS
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/En_clk_din/En_clk_din.sym # of pins=7
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/En_clk_din/En_clk_din.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/En_clk_din/En_clk_din.sch
.subckt En_clk_din VDD VSS clk clock enable D_in Data_in
*.PININFO D_in:I enable:I clk:B VDD:B VSS:B clock:O Data_in:O
x6 net1 D_in Data_in VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__and2_1
x15 enable net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x2 net2 clk clock VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__and2_1
x3 enable net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
* noconn VSS
* noconn VDD
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_not/not.sym # of pins=4
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_not/not.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_not/not.sch
.subckt not vdd in out vss
*.PININFO vdd:B vss:B in:B out:B
XM1 out in vdd vdd pfet_03v3 L=0.35u W=1u nf=1 m=1
XM3 out in vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_nor/nor.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_nor/nor.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_nor/nor.sch
.subckt nor vdd vss A B Z
*.PININFO vdd:B vss:B A:I Z:O B:I
XM1 net1 A vdd vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
XM3 Z B vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM2 Z A vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM4 Z B net1 vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_monostable/monostable.sym # of pins=7
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_monostable/monostable.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_monostable/monostable.sch
.subckt monostable vss vdd vin vres phi_1 phi_2 vneg
*.PININFO vin:I vdd:B vss:B phi_1:O vres:I phi_2:O vneg:O
x2 vdd net2 vneg vss not
XM2 net2 vres vss vss nfet_03v3 L=0.3u W=1u nf=1 m=1
x13 vdd vss net1 vneg vin nand
x14 vdd vneg phi_1 vss not
XC2 net1 net2 cap_mim_2f0fF c_width=5e-6 c_length=5e-6 m=1
x1 vdd net5 net3 vss not
XM1 net5 vres vss vss nfet_03v3 L=0.3u W=1u nf=1 m=1
x3 vdd vss net4 net3 phi_1 nand
x4 vdd net3 phi_2 vss not
XC1 net4 net5 cap_mim_2f0fF c_width=5e-6 c_length=5e-6 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_refractory/refractory.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_refractory/refractory.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_refractory/refractory.sch
.subckt refractory vss vdd vspike_down vneg vrefrac
*.PININFO vspike_down:I vdd:B vss:B vrefrac:O vneg:I
x22 vdd vrefrac net2 net1 vss ota_1stage
XM9 net1 net1 vrefrac vss nfet_03v3 L=0.5u W=0.5u nf=1 m=1
XM10 vspike_down vspike_down net1 vss nfet_03v3 L=0.5u W=0.5u nf=1 m=1
XM11 vneg vneg net2 vss nfet_03v3 L=13u W=0.36u nf=1 m=1
XM12 net2 net2 vss vss nfet_03v3 L=0.28u W=15u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_vdiv/nvdiv.sym # of pins=6
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_vdiv/nvdiv.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_vdiv/nvdiv.sch
.subckt nvdiv vss vdd vref vspike_up vspike_down vres
*.PININFO vref:O vdd:B vss:B vspike_up:O vspike_down:O vres:O
XM15 vdd vdd vspike_up vss nfet_03v3 L=0.28u W=0.36u nf=1 m=1
XM18 vspike_down vspike_down vres vss nfet_03v3 L=0.5u W=0.5u nf=1 m=1
XM16 vp vp vspike_down vss nfet_03v3 L=0.5u W=0.5u nf=1 m=1
XM19 vres vres vss vss nfet_03v3 L=0.8u W=0.5u nf=1 m=1
XM17 vspike_up vspike_up vp vss nfet_03v3 L=0.28u W=0.36u nf=1 m=1
XM20 vref vref vss vss nfet_03v3 L=0.28u W=0.36u nf=1 m=1
XM21 vdd vdd vref vss nfet_03v3 L=0.28u W=0.55u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sch
.subckt ShiftReg_row_10_2 D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8]
+ gc[9] gc[10] PHI_1 PHI_2 EN VDD VSS
*.PININFO PHI_1:I PHI_2:I D_in:I Q[1:10]:O VDD:B VSS:B EN:B gc[1:10]:B
xFF[1] Q[1] D_in PHI_1 gc[1] PHI_2 EN VDD VSS DFF_2phase_1
xFF[2] Q[2] Q[1] PHI_1 gc[2] PHI_2 EN VDD VSS DFF_2phase_1
xFF[3] Q[3] Q[2] PHI_1 gc[3] PHI_2 EN VDD VSS DFF_2phase_1
xFF[4] Q[4] Q[3] PHI_1 gc[4] PHI_2 EN VDD VSS DFF_2phase_1
xFF[5] Q[5] Q[4] PHI_1 gc[5] PHI_2 EN VDD VSS DFF_2phase_1
xFF[6] Q[6] Q[5] PHI_1 gc[6] PHI_2 EN VDD VSS DFF_2phase_1
xFF[7] Q[7] Q[6] PHI_1 gc[7] PHI_2 EN VDD VSS DFF_2phase_1
xFF[8] Q[8] Q[7] PHI_1 gc[8] PHI_2 EN VDD VSS DFF_2phase_1
xFF[9] Q[9] Q[8] PHI_1 gc[9] PHI_2 EN VDD VSS DFF_2phase_1
xFF[10] Q[10] Q[9] PHI_1 gc[10] PHI_2 EN VDD VSS DFF_2phase_1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sch
.subckt swmatrix_Tgate gated_control T2 T1 VSS VDD
*.PININFO T1:B T2:B VDD:B VSS:B gated_control:I
XM1 T1 gated_control T2 VSS nfet_03v3 L=0.28u W=24u nf=6 m=1
XM2 T1 gated_controlb T2 VDD pfet_03v3 L=0.28u W=72u nf=6 m=1
**** begin user architecture code
**** end user architecture code
x1 gated_control gated_controlb VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends


* expanding   symbol:  designs/libs/core_LIF_comp/core_nand/nand.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_nand/nand.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/core_LIF_comp/core_nand/nand.sch
.subckt nand vdd vss Z A B
*.PININFO vdd:B vss:B A:I Z:O B:I
XM1 Z A vdd vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
XM3 net1 B vss vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM2 Z A net1 vss nfet_03v3 L=0.28u W=1u nf=1 m=1
XM4 Z B vdd vdd pfet_03v3 L=0.28u W=1u nf=1 m=1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 Q D PHI_1 gated_control PHI_2 EN VDD VSS
*.PININFO D:I PHI_1:I PHI_2:I Q:O VDD:B VSS:B gated_control:O EN:I
xmain D PHI_1 out_m VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
* noconn VSS
* noconn VDD
x1 net1 gated_control VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x2 EN Q net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
.ends

