magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
rect 0 0 3 2
<< l34d0 >>
<< l36d0 >>
<< l42d0 >>
<< l46d0 >>
<< l81d0 >>
<< labels >>
rlabel l34d10 2.149 1.112 2.149 1.112 0 vss
rlabel l34d10 2.1425 1.6295 2.1425 1.6295 0 vdd
rlabel l34d10 0.62 1.34 0.62 1.34 0 vin
rlabel l34d10 2.7815 1.315 2.7815 1.315 0 phi_2
rlabel l34d10 1.372 0.792 1.372 0.792 0 vres
rlabel l34d10 2.6045 0.793 2.6045 0.793 0 vres
rlabel l36d10 0.9765 1.396 0.9765 1.396 0 vneg
rlabel l36d10 1.638 1.3105 1.638 1.3105 0 phi_1
use nand nand_1
timestamp 1757365861
transform -1 0 1 0 1 2
box 0 0 0 0
use not not_1
timestamp 1757365861
transform -1 0 1 0 1 2
box 0 0 0 0
use not not_2
timestamp 1757365861
transform -1 0 1 0 1 2
box 0 0 0 0
use via_devx2418 via_devx2418_1
timestamp 1757365861
transform 1 0 0 0 1 1
box 0 0 0 0
use via_devx2419 via_devx2419_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2419 via_devx2419_2
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2420 via_devx2420_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2418 via_devx2418_2
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use cap_mim cap_mim_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 1 1
use via_devx2421 via_devx2421_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2422 via_devx2422_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2423 via_devx2423_1
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use nand nand_2
timestamp 1757365861
transform -1 0 2 0 1 2
box 0 0 0 0
use not not_3
timestamp 1757365861
transform -1 0 2 0 1 2
box 0 0 0 0
use not not_4
timestamp 1757365861
transform -1 0 3 0 1 2
box 0 0 0 0
use via_devx2424 via_devx2424_1
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_1
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2420 via_devx2420_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2424 via_devx2424_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use cap_mim cap_mim_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 1 1
use via_devx2421 via_devx2421_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2422 via_devx2422_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2424 via_devx2424_3
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_2
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_3
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
use via_devx2420 via_devx2420_3
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use nfetx2415 nfetx2415_1
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2420 via_devx2420_4
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use nfetx2415 nfetx2415_2
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_4
timestamp 1757365861
transform 1 0 1 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_5
timestamp 1757365861
transform 1 0 3 0 1 1
box 0 0 0 0
use via_devx2425 via_devx2425_6
timestamp 1757365861
transform 1 0 2 0 1 1
box 0 0 0 0
<< end >>
