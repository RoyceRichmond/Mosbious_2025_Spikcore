magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l34d0 >>
<< l21d0 >>
<< l36d0 >>
<< labels >>
rlabel l34d10 0.016 -0.1735 0.016 -0.1735 0 A
rlabel l34d10 0.125 -0.176 0.125 -0.176 0 B
rlabel l34d10 -0.104 -0.1815 -0.104 -0.1815 0 Z
rlabel l34d10 0.102 -0.4185 0.102 -0.4185 0 vss
rlabel l34d10 0.094 0.107 0.094 0.107 0 vdd
use pfetx246 pfetx246_1
timestamp 1757365861
transform 1 0 1 0 1 0
box 0 0 0 0
use pfetx247 pfetx247_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2415 via_devx2415_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use pfetx248 pfetx248_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2416 via_devx2416_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2416 via_devx2416_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2412 nfetx2412_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2416 via_devx2416_3
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2413 nfetx2413_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2416 via_devx2416_4
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
<< end >>
