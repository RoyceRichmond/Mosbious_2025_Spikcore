* NGSPICE file created from TG_bootstrapped.ext - technology: gf180mcuD

.subckt TG_bootstrapped_pex vdd vss clk nclk vin vout
X0 vout.t35 a_5673_n171.t4 vin.t29 vss.t27 nfet_03v3 ad=2.38815p pd=9.05u as=1.0179p ps=4.435u w=3.915u l=0.42u
X1 vin.t35 a_5673_n171.t5 vout.t34 vss.t26 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X2 vin.t3 a_5297_1329.t4 vout.t1 vdd.t25 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X3 a_8039_2775# a_5944_2887# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X4 vin.t8 clk.t0 a_8039_2775# vss.t9 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X5 vin.t5 a_5297_1329.t5 vout.t3 vdd.t24 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X6 vout.t2 a_5297_1329.t6 vin.t4 vdd.t23 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X7 vout.t0 a_5297_1329.t7 vin.t0 vdd.t22 pfet_03v3 ad=2.028p pd=7.54u as=0.8112p ps=3.64u w=3.12u l=0.42u
X8 vin.t6 a_5297_1329.t8 vout.t4 vdd.t21 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X9 vin.t23 a_5297_1329.t9 vout.t19 vdd.t20 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X10 vss.t4 nclk.t0 a_5673_n171.t1 vss.t3 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X11 vout.t18 a_5297_1329.t10 vin.t22 vdd.t19 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X12 vin.t21 a_5297_1329.t11 vout.t17 vdd.t18 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X13 vin.t13 a_5297_1329.t12 vout.t9 vdd.t17 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X14 a_8034_n1134# nclk.t1 vss.t2 vss.t1 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X15 vin.t1 nclk.t2 a_8034_n1134# vdd.t1 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X16 vin.t32 a_5673_n171.t6 vout.t33 vss.t25 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X17 vout.t32 a_5673_n171.t7 vin.t37 vss.t24 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X18 vout.t31 a_5673_n171.t8 vin.t31 vss.t23 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X19 vout.t30 a_5673_n171.t9 vin.t27 vss.t22 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X20 vdd.t28 clk.t1 a_5297_1329.t3 vdd.t27 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X21 vin.t36 a_5673_n171.t10 vout.t29 vss.t21 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X22 a_5904_n1280# clk.t2 vss.t8 vss.t7 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X23 a_5297_1329.t1 nclk.t3 a_5944_2887# vdd.t5 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X24 a_5673_n171.t0 nclk.t4 a_5904_n1280# vdd.t26 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X25 vin.t20 a_5297_1329.t13 vout.t16 vdd.t16 pfet_03v3 ad=0.8112p pd=3.64u as=2.028p ps=7.54u w=3.12u l=0.42u
X26 vout.t10 a_5297_1329.t14 vin.t14 vdd.t15 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X27 vout.t15 a_5297_1329.t15 vin.t19 vdd.t14 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X28 vout.t8 a_5297_1329.t16 vin.t12 vdd.t13 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X29 vin.t18 a_5297_1329.t17 vout.t14 vdd.t12 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X30 a_8034_n1134# a_5904_n1280# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X31 vin.t2 nclk.t5 a_8039_2775# vdd.t2 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X32 vdd.t0 nclk.t6 a_5297_1329.t0 vss.t0 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X33 a_5297_1329.t2 clk.t3 a_5944_2887# vss.t6 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X34 vin.t24 a_5673_n171.t11 vout.t28 vss.t20 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X35 vss.t10 clk.t4 a_5673_n171.t2 vdd.t29 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X36 vin.t28 a_5673_n171.t12 vout.t27 vss.t19 nfet_03v3 ad=1.0179p pd=4.435u as=2.38815p ps=9.05u w=3.915u l=0.42u
X37 vin.t38 a_5673_n171.t13 vout.t26 vss.t18 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X38 vout.t25 a_5673_n171.t14 vin.t25 vss.t17 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X39 vdd.t4 nclk.t7 a_8039_2775# vdd.t3 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X40 vout.t24 a_5673_n171.t15 vin.t39 vss.t16 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X41 vout.t7 a_5297_1329.t18 vin.t11 vdd.t11 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X42 vin.t17 a_5297_1329.t19 vout.t13 vdd.t10 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X43 a_5944_2887# clk.t5 vdd.t31 vdd.t30 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X44 vout.t5 a_5297_1329.t20 vin.t9 vdd.t9 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X45 vout.t12 a_5297_1329.t21 vin.t16 vdd.t8 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X46 vout.t6 a_5297_1329.t22 vin.t10 vdd.t7 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X47 vin.t15 a_5297_1329.t23 vout.t11 vdd.t6 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X48 vout.t23 a_5673_n171.t16 vin.t30 vss.t15 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X49 vin.t7 clk.t6 a_8034_n1134# vss.t5 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X50 vout.t22 a_5673_n171.t17 vin.t34 vss.t14 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X51 vin.t26 a_5673_n171.t18 vout.t21 vss.t13 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X52 vin.t33 a_5673_n171.t19 vout.t20 vss.t12 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X53 a_5673_n171.t3 clk.t7 a_5904_n1280# vss.t11 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
R0 a_5673_n171.n5 a_5673_n171.t12 50.5346
R1 a_5673_n171.n14 a_5673_n171.t4 50.5346
R2 a_5673_n171.n5 a_5673_n171.t17 50.3231
R3 a_5673_n171.n6 a_5673_n171.t5 50.3231
R4 a_5673_n171.n7 a_5673_n171.t8 50.3231
R5 a_5673_n171.n8 a_5673_n171.t13 50.3231
R6 a_5673_n171.n9 a_5673_n171.t16 50.3231
R7 a_5673_n171.n12 a_5673_n171.t6 50.3231
R8 a_5673_n171.n11 a_5673_n171.t9 50.3231
R9 a_5673_n171.n20 a_5673_n171.t10 50.3231
R10 a_5673_n171.n19 a_5673_n171.t15 50.3231
R11 a_5673_n171.n18 a_5673_n171.t18 50.3231
R12 a_5673_n171.n17 a_5673_n171.t7 50.3231
R13 a_5673_n171.n16 a_5673_n171.t11 50.3231
R14 a_5673_n171.n15 a_5673_n171.t14 50.3231
R15 a_5673_n171.n14 a_5673_n171.t19 50.3231
R16 a_5673_n171.n28 a_5673_n171.t3 9.65132
R17 a_5673_n171.n3 a_5673_n171.t1 9.65118
R18 a_5673_n171.n22 a_5673_n171.n10 9.0005
R19 a_5673_n171.n22 a_5673_n171.n13 9.0005
R20 a_5673_n171.n22 a_5673_n171.n4 9.0005
R21 a_5673_n171.n22 a_5673_n171.n21 9.0005
R22 a_5673_n171.n25 a_5673_n171.n23 4.5005
R23 a_5673_n171.n26 a_5673_n171.n2 4.5005
R24 a_5673_n171.n27 a_5673_n171.n26 4.5005
R25 a_5673_n171.n26 a_5673_n171.n25 4.5005
R26 a_5673_n171.n3 a_5673_n171.t2 3.70851
R27 a_5673_n171.t0 a_5673_n171.n28 3.70835
R28 a_5673_n171.n24 a_5673_n171.n1 2.24455
R29 a_5673_n171.n23 a_5673_n171.n0 2.24204
R30 a_5673_n171.n25 a_5673_n171.n3 1.04078
R31 a_5673_n171.n28 a_5673_n171.n27 1.03838
R32 a_5673_n171.n15 a_5673_n171.n14 0.212
R33 a_5673_n171.n16 a_5673_n171.n15 0.212
R34 a_5673_n171.n17 a_5673_n171.n16 0.212
R35 a_5673_n171.n18 a_5673_n171.n17 0.212
R36 a_5673_n171.n19 a_5673_n171.n18 0.212
R37 a_5673_n171.n9 a_5673_n171.n8 0.212
R38 a_5673_n171.n8 a_5673_n171.n7 0.212
R39 a_5673_n171.n7 a_5673_n171.n6 0.212
R40 a_5673_n171.n6 a_5673_n171.n5 0.212
R41 a_5673_n171.n21 a_5673_n171.n20 0.147875
R42 a_5673_n171.n11 a_5673_n171.n4 0.134375
R43 a_5673_n171.n23 a_5673_n171.n22 0.122181
R44 a_5673_n171.n13 a_5673_n171.n12 0.120875
R45 a_5673_n171.n10 a_5673_n171.n9 0.107375
R46 a_5673_n171.n12 a_5673_n171.n10 0.105125
R47 a_5673_n171.n13 a_5673_n171.n11 0.091625
R48 a_5673_n171.n20 a_5673_n171.n4 0.078125
R49 a_5673_n171.n21 a_5673_n171.n19 0.064625
R50 a_5673_n171.n25 a_5673_n171.n24 0.0365
R51 a_5673_n171.n24 a_5673_n171.n2 0.0365
R52 a_5673_n171.n27 a_5673_n171.n0 0.0189283
R53 a_5673_n171.n2 a_5673_n171.n0 0.0189283
R54 a_5673_n171.n26 a_5673_n171.n1 0.013894
R55 a_5673_n171.n23 a_5673_n171.n1 0.013894
R56 vin.n80 vin.t8 13.8016
R57 vin.n87 vin.t7 9.92542
R58 vin vin.n86 9.75035
R59 vin.n81 vin.n80 4.99212
R60 vin.n83 vin.n82 4.60986
R61 vin.n84 vin.n83 4.5696
R62 vin.n85 vin.n84 4.5005
R63 vin.n82 vin.n81 4.5005
R64 vin.n83 vin.t2 3.48383
R65 vin.n87 vin.t1 3.48383
R66 vin.n5 vin.n3 2.12064
R67 vin.n46 vin.n44 2.12064
R68 vin.n5 vin.n4 2.05296
R69 vin.n76 vin.n75 2.05296
R70 vin.n69 vin.n68 2.05296
R71 vin.n15 vin.n14 2.05296
R72 vin.n61 vin.n60 2.05296
R73 vin.n35 vin.n34 2.05296
R74 vin.n53 vin.n52 2.05296
R75 vin.n46 vin.n45 2.05296
R76 vin.n1 vin.n0 1.87421
R77 vin.n43 vin.n42 1.86774
R78 vin.n9 vin.n8 1.86521
R79 vin.n17 vin.n16 1.86521
R80 vin.n21 vin.n20 1.86521
R81 vin.n27 vin.n26 1.86521
R82 vin.n31 vin.n30 1.86521
R83 vin.n39 vin.n38 1.86521
R84 vin.n48 vin.n47 1.5005
R85 vin.n49 vin.n36 1.5005
R86 vin.n51 vin.n50 1.5005
R87 vin.n54 vin.n33 1.5005
R88 vin.n56 vin.n55 1.5005
R89 vin.n57 vin.n24 1.5005
R90 vin.n59 vin.n58 1.5005
R91 vin.n62 vin.n23 1.5005
R92 vin.n64 vin.n63 1.5005
R93 vin.n66 vin.n65 1.5005
R94 vin.n67 vin.n13 1.5005
R95 vin.n71 vin.n70 1.5005
R96 vin.n72 vin.n6 1.5005
R97 vin.n74 vin.n73 1.5005
R98 vin.n77 vin.n2 1.5005
R99 vin.n79 vin.n78 1.5005
R100 vin.n48 vin.n43 1.1255
R101 vin.n49 vin.n41 1.1255
R102 vin.n50 vin.n40 1.1255
R103 vin.n37 vin.n33 1.1255
R104 vin.n56 vin.n32 1.1255
R105 vin.n57 vin.n29 1.1255
R106 vin.n58 vin.n28 1.1255
R107 vin.n25 vin.n23 1.1255
R108 vin.n64 vin.n22 1.1255
R109 vin.n65 vin.n19 1.1255
R110 vin.n18 vin.n13 1.1255
R111 vin.n71 vin.n12 1.1255
R112 vin.n72 vin.n11 1.1255
R113 vin.n73 vin.n10 1.1255
R114 vin.n7 vin.n2 1.1255
R115 vin.n79 vin.n1 1.1255
R116 vin.n86 vin.n85 1.04563
R117 vin.n48 vin 0.601237
R118 vin.n44 vin.t9 0.583833
R119 vin.n44 vin.t20 0.583833
R120 vin.n45 vin.t14 0.583833
R121 vin.n45 vin.t5 0.583833
R122 vin.n52 vin.t22 0.583833
R123 vin.n52 vin.t15 0.583833
R124 vin.n34 vin.t16 0.583833
R125 vin.n34 vin.t18 0.583833
R126 vin.n60 vin.t19 0.583833
R127 vin.n60 vin.t6 0.583833
R128 vin.n14 vin.t12 0.583833
R129 vin.n14 vin.t23 0.583833
R130 vin.n68 vin.t4 0.583833
R131 vin.n68 vin.t17 0.583833
R132 vin.n75 vin.t10 0.583833
R133 vin.n75 vin.t21 0.583833
R134 vin.n4 vin.t11 0.583833
R135 vin.n4 vin.t13 0.583833
R136 vin.n3 vin.t0 0.583833
R137 vin.n3 vin.t3 0.583833
R138 vin.n42 vin.t34 0.418891
R139 vin.n42 vin.t28 0.418891
R140 vin.n38 vin.t31 0.418891
R141 vin.n38 vin.t35 0.418891
R142 vin.n30 vin.t30 0.418891
R143 vin.n30 vin.t38 0.418891
R144 vin.n26 vin.t27 0.418891
R145 vin.n26 vin.t32 0.418891
R146 vin.n20 vin.t39 0.418891
R147 vin.n20 vin.t36 0.418891
R148 vin.n16 vin.t37 0.418891
R149 vin.n16 vin.t26 0.418891
R150 vin.n8 vin.t25 0.418891
R151 vin.n8 vin.t24 0.418891
R152 vin.n0 vin.t29 0.418891
R153 vin.n0 vin.t33 0.418891
R154 vin vin.n87 0.394842
R155 vin.n85 vin.n81 0.1805
R156 vin.n84 vin 0.096125
R157 vin.n82 vin 0.084875
R158 vin.n80 vin 0.037625
R159 vin.n78 vin.n77 0.0311
R160 vin.n74 vin.n6 0.0311
R161 vin.n70 vin.n6 0.0311
R162 vin.n67 vin.n66 0.0311
R163 vin.n63 vin.n62 0.0311
R164 vin.n59 vin.n24 0.0311
R165 vin.n55 vin.n54 0.0311
R166 vin.n51 vin.n36 0.0311
R167 vin.n47 vin.n36 0.0311
R168 vin.n69 vin.n67 0.02966
R169 vin.n54 vin.n53 0.02786
R170 vin.n77 vin.n76 0.02606
R171 vin.n7 vin.n1 0.0244062
R172 vin.n11 vin.n10 0.0244062
R173 vin.n12 vin.n11 0.0244062
R174 vin.n19 vin.n18 0.0244062
R175 vin.n25 vin.n22 0.0244062
R176 vin.n29 vin.n28 0.0244062
R177 vin.n37 vin.n32 0.0244062
R178 vin.n41 vin.n40 0.0244062
R179 vin.n43 vin.n41 0.0244062
R180 vin.n18 vin.n17 0.0232812
R181 vin.n63 vin.n15 0.02318
R182 vin.n39 vin.n37 0.021875
R183 vin.n35 vin.n24 0.02138
R184 vin.n9 vin.n7 0.0204687
R185 vin.n22 vin.n21 0.0182187
R186 vin.n31 vin.n29 0.0168125
R187 vin.n61 vin.n59 0.0167
R188 vin.n62 vin.n61 0.0149
R189 vin.n28 vin.n27 0.0131563
R190 vin.n78 vin.n5 0.01202
R191 vin.n27 vin.n25 0.01175
R192 vin.n55 vin.n35 0.01022
R193 vin.n79 vin.n2 0.0084729
R194 vin.n73 vin.n2 0.0084729
R195 vin.n73 vin.n72 0.0084729
R196 vin.n72 vin.n71 0.0084729
R197 vin.n71 vin.n13 0.0084729
R198 vin.n65 vin.n13 0.0084729
R199 vin.n65 vin.n64 0.0084729
R200 vin.n64 vin.n23 0.0084729
R201 vin.n58 vin.n23 0.0084729
R202 vin.n58 vin.n57 0.0084729
R203 vin.n57 vin.n56 0.0084729
R204 vin.n56 vin.n33 0.0084729
R205 vin.n50 vin.n33 0.0084729
R206 vin.n50 vin.n49 0.0084729
R207 vin.n49 vin.n48 0.0084729
R208 vin.n66 vin.n15 0.00842
R209 vin.n32 vin.n31 0.00809375
R210 vin.n21 vin.n19 0.0066875
R211 vin.n76 vin.n74 0.00554
R212 vin.n10 vin.n9 0.0044375
R213 vin.n53 vin.n51 0.00374
R214 vin.n47 vin.n46 0.00374
R215 vin.n40 vin.n39 0.00303125
R216 vin.n86 vin.n79 0.00218838
R217 vin.n70 vin.n69 0.00194
R218 vin.n17 vin.n12 0.001625
R219 vout.n1 vout.t0 2.56303
R220 vout.n28 vout.t16 2.56303
R221 vout.n29 vout.n26 2.31025
R222 vout.n31 vout.n26 2.2505
R223 vout.n33 vout.n32 2.2505
R224 vout.n35 vout.n34 2.2505
R225 vout.n36 vout.n20 2.2505
R226 vout.n39 vout.n38 2.2505
R227 vout.n40 vout.n19 2.2505
R228 vout.n42 vout.n41 2.2505
R229 vout.n44 vout.n16 2.2505
R230 vout.n46 vout.n45 2.2505
R231 vout.n48 vout.n47 2.2505
R232 vout.n49 vout.n10 2.2505
R233 vout.n52 vout.n51 2.2505
R234 vout.n53 vout.n9 2.2505
R235 vout.n55 vout.n54 2.2505
R236 vout.n57 vout.n6 2.2505
R237 vout.n59 vout.n58 2.2505
R238 vout.n61 vout.n60 2.2505
R239 vout.n62 vout.n0 2.2505
R240 vout.n65 vout.n64 2.2505
R241 vout.n28 vout.t27 2.24523
R242 vout.n1 vout.t35 2.24523
R243 vout.n5 vout.n4 1.60155
R244 vout.n56 vout.n8 1.60155
R245 vout.n50 vout.n12 1.60155
R246 vout.n15 vout.n14 1.60155
R247 vout.n43 vout.n18 1.60155
R248 vout.n37 vout.n22 1.60155
R249 vout.n25 vout.n24 1.60155
R250 vout.n63 vout.n2 1.47822
R251 vout.n5 vout.n3 1.47822
R252 vout.n56 vout.n7 1.47822
R253 vout.n50 vout.n11 1.47822
R254 vout.n15 vout.n13 1.47822
R255 vout.n43 vout.n17 1.47822
R256 vout.n37 vout.n21 1.47822
R257 vout.n25 vout.n23 1.47822
R258 vout.n30 vout.n27 1.47822
R259 vout vout.n65 1.02411
R260 vout.n2 vout.t1 0.583833
R261 vout.n2 vout.t7 0.583833
R262 vout.n3 vout.t9 0.583833
R263 vout.n3 vout.t6 0.583833
R264 vout.n7 vout.t17 0.583833
R265 vout.n7 vout.t2 0.583833
R266 vout.n11 vout.t13 0.583833
R267 vout.n11 vout.t8 0.583833
R268 vout.n13 vout.t19 0.583833
R269 vout.n13 vout.t15 0.583833
R270 vout.n17 vout.t4 0.583833
R271 vout.n17 vout.t12 0.583833
R272 vout.n21 vout.t14 0.583833
R273 vout.n21 vout.t18 0.583833
R274 vout.n23 vout.t11 0.583833
R275 vout.n23 vout.t10 0.583833
R276 vout.n27 vout.t3 0.583833
R277 vout.n27 vout.t5 0.583833
R278 vout.n4 vout.t20 0.418891
R279 vout.n4 vout.t25 0.418891
R280 vout.n8 vout.t28 0.418891
R281 vout.n8 vout.t32 0.418891
R282 vout.n12 vout.t21 0.418891
R283 vout.n12 vout.t24 0.418891
R284 vout.n14 vout.t29 0.418891
R285 vout.n14 vout.t30 0.418891
R286 vout.n18 vout.t33 0.418891
R287 vout.n18 vout.t23 0.418891
R288 vout.n22 vout.t26 0.418891
R289 vout.n22 vout.t31 0.418891
R290 vout.n24 vout.t34 0.418891
R291 vout.n24 vout.t22 0.418891
R292 vout.n62 vout.n61 0.0605
R293 vout.n58 vout.n57 0.0605
R294 vout.n55 vout.n9 0.0605
R295 vout.n51 vout.n9 0.0605
R296 vout.n49 vout.n48 0.0605
R297 vout.n45 vout.n44 0.0605
R298 vout.n42 vout.n19 0.0605
R299 vout.n38 vout.n19 0.0605
R300 vout.n36 vout.n35 0.0605
R301 vout.n32 vout.n31 0.0605
R302 vout.n65 vout.n0 0.060251
R303 vout.n60 vout.n0 0.060251
R304 vout.n60 vout.n59 0.060251
R305 vout.n59 vout.n6 0.060251
R306 vout.n54 vout.n6 0.060251
R307 vout.n54 vout.n53 0.060251
R308 vout.n53 vout.n52 0.060251
R309 vout.n52 vout.n10 0.060251
R310 vout.n47 vout.n10 0.060251
R311 vout.n47 vout.n46 0.060251
R312 vout.n46 vout.n16 0.060251
R313 vout.n41 vout.n16 0.060251
R314 vout.n41 vout.n40 0.060251
R315 vout.n40 vout.n39 0.060251
R316 vout.n39 vout.n20 0.060251
R317 vout.n34 vout.n20 0.060251
R318 vout.n34 vout.n33 0.060251
R319 vout.n33 vout.n26 0.060251
R320 vout.n63 vout.n62 0.05525
R321 vout.n31 vout.n30 0.05375
R322 vout.n50 vout.n49 0.05225
R323 vout.n44 vout.n43 0.05075
R324 vout.n37 vout.n36 0.04925
R325 vout.n57 vout.n56 0.04775
R326 vout.n58 vout.n5 0.03425
R327 vout.n35 vout.n25 0.03275
R328 vout.n45 vout.n15 0.03125
R329 vout.n48 vout.n15 0.02975
R330 vout.n32 vout.n25 0.02825
R331 vout.n61 vout.n5 0.02675
R332 vout.n56 vout.n55 0.01325
R333 vout.n38 vout.n37 0.01175
R334 vout.n43 vout.n42 0.01025
R335 vout.n51 vout.n50 0.00875
R336 vout.n30 vout.n29 0.00725
R337 vout.n64 vout.n1 0.00575
R338 vout.n64 vout.n63 0.00575
R339 vout.n29 vout.n28 0.00425
R340 vss.n14 vss.n13 28130.3
R341 vss.n13 vss.n3 3658.85
R342 vss.n15 vss.n14 3473.68
R343 vss.n14 vss.t6 2794.63
R344 vss.n13 vss.t1 2578.99
R345 vss.t5 vss.t3 1060.25
R346 vss.t9 vss.t0 920.038
R347 vss.n12 vss.t11 541.668
R348 vss.t3 vss.n20 480.928
R349 vss.n20 vss.t11 480.928
R350 vss.n23 vss.t5 470.882
R351 vss.t0 vss.n2 416.243
R352 vss.t6 vss.n2 416.243
R353 vss.n3 vss.t9 406.25
R354 vss.n24 vss.t27 358.844
R355 vss.t12 vss.t27 319.728
R356 vss.t17 vss.t12 319.728
R357 vss.t20 vss.t17 319.728
R358 vss.t24 vss.t20 319.728
R359 vss.t13 vss.t24 319.728
R360 vss.t16 vss.t13 319.728
R361 vss.t21 vss.t16 319.728
R362 vss.t22 vss.t21 319.728
R363 vss.t25 vss.t22 319.728
R364 vss.t15 vss.t25 319.728
R365 vss.t18 vss.t15 319.728
R366 vss.t23 vss.t18 319.728
R367 vss.n24 vss.n23 301.611
R368 vss.t1 vss.n7 175.298
R369 vss.t14 vss.t26 131.823
R370 vss.n12 vss.t23 122.45
R371 vss.t19 vss.t7 112.891
R372 vss.n25 vss.n7 86.9476
R373 vss.t26 vss.n12 81.3381
R374 vss.n15 vss.t19 62.4061
R375 vss.n25 vss.n24 37.1634
R376 vss.n28 vss.n3 19.8888
R377 vss.n23 vss.n22 19.6851
R378 vss.t7 vss.t14 18.9325
R379 vss.n17 vss.n16 11.0839
R380 vss.n16 vss.t8 10.8815
R381 vss.n21 vss.t2 10.877
R382 vss.n21 vss.n7 10.4837
R383 vss.n16 vss.n15 10.4793
R384 vss.n5 vss.t4 9.6559
R385 vss.n22 vss.n21 9.22213
R386 vss.n33 vss.n32 4.59325
R387 vss.n10 vss.n8 4.59325
R388 vss.n31 vss.n30 4.5005
R389 vss.n19 vss.n18 4.5005
R390 vss.n11 vss.n9 4.5005
R391 vss.n18 vss.n17 4.5005
R392 vss.n1 vss.n0 4.5005
R393 vss.n30 vss.n29 4.5005
R394 vss.n26 vss.n25 3.80854
R395 vss.n5 vss.t10 3.71674
R396 vss.n6 vss.n5 2.94978
R397 vss.n32 vss.n31 2.20487
R398 vss.n19 vss.n8 2.20487
R399 vss.n26 vss.n6 1.34213
R400 vss.n27 vss.n4 1.02307
R401 vss.n28 vss.n27 0.918196
R402 vss vss.n33 0.60333
R403 vss.n22 vss.n4 0.4415
R404 vss.n31 vss.n2 0.298561
R405 vss.n29 vss.n28 0.280052
R406 vss.n20 vss.n19 0.271533
R407 vss.n27 vss.n26 0.201851
R408 vss.n30 vss.n1 0.188872
R409 vss.n18 vss.n9 0.188872
R410 vss.n22 vss.n6 0.176
R411 vss.n10 vss.n4 0.0973229
R412 vss.n32 vss.n1 0.0932551
R413 vss.n9 vss.n8 0.0932551
R414 vss.n29 vss.n0 0.0387075
R415 vss.n33 vss.n0 0.0387075
R416 vss.n11 vss.n10 0.0116647
R417 vss.n17 vss.n11 0.0116647
R418 a_5297_1329.n6 a_5297_1329.t13 43.8541
R419 a_5297_1329.n17 a_5297_1329.t7 43.8541
R420 a_5297_1329.n6 a_5297_1329.t20 43.6315
R421 a_5297_1329.n7 a_5297_1329.t5 43.6315
R422 a_5297_1329.n8 a_5297_1329.t14 43.6315
R423 a_5297_1329.n9 a_5297_1329.t23 43.6315
R424 a_5297_1329.n10 a_5297_1329.t10 43.6315
R425 a_5297_1329.n11 a_5297_1329.t17 43.6315
R426 a_5297_1329.n12 a_5297_1329.t21 43.6315
R427 a_5297_1329.n15 a_5297_1329.t8 43.6315
R428 a_5297_1329.n14 a_5297_1329.t15 43.6315
R429 a_5297_1329.n25 a_5297_1329.t9 43.6315
R430 a_5297_1329.n24 a_5297_1329.t16 43.6315
R431 a_5297_1329.n23 a_5297_1329.t19 43.6315
R432 a_5297_1329.n22 a_5297_1329.t6 43.6315
R433 a_5297_1329.n21 a_5297_1329.t11 43.6315
R434 a_5297_1329.n20 a_5297_1329.t22 43.6315
R435 a_5297_1329.n19 a_5297_1329.t12 43.6315
R436 a_5297_1329.n18 a_5297_1329.t18 43.6315
R437 a_5297_1329.n17 a_5297_1329.t4 43.6315
R438 a_5297_1329.n3 a_5297_1329.t2 9.65161
R439 a_5297_1329.t0 a_5297_1329.n32 9.65118
R440 a_5297_1329.n27 a_5297_1329.n13 9.0005
R441 a_5297_1329.n27 a_5297_1329.n16 9.0005
R442 a_5297_1329.n27 a_5297_1329.n5 9.0005
R443 a_5297_1329.n27 a_5297_1329.n26 9.0005
R444 a_5297_1329.n31 a_5297_1329.n0 4.5005
R445 a_5297_1329.n30 a_5297_1329.n29 4.5005
R446 a_5297_1329.n30 a_5297_1329.n4 4.5005
R447 a_5297_1329.n31 a_5297_1329.n30 4.5005
R448 a_5297_1329.n32 a_5297_1329.t3 3.70851
R449 a_5297_1329.n3 a_5297_1329.t1 3.7081
R450 a_5297_1329.n2 a_5297_1329.n1 2.24497
R451 a_5297_1329.n28 a_5297_1329.n0 2.24204
R452 a_5297_1329.n32 a_5297_1329.n31 1.04078
R453 a_5297_1329.n4 a_5297_1329.n3 1.03844
R454 a_5297_1329.n12 a_5297_1329.n11 0.223132
R455 a_5297_1329.n11 a_5297_1329.n10 0.223132
R456 a_5297_1329.n10 a_5297_1329.n9 0.223132
R457 a_5297_1329.n9 a_5297_1329.n8 0.223132
R458 a_5297_1329.n8 a_5297_1329.n7 0.223132
R459 a_5297_1329.n7 a_5297_1329.n6 0.223132
R460 a_5297_1329.n18 a_5297_1329.n17 0.223132
R461 a_5297_1329.n19 a_5297_1329.n18 0.223132
R462 a_5297_1329.n20 a_5297_1329.n19 0.223132
R463 a_5297_1329.n21 a_5297_1329.n20 0.223132
R464 a_5297_1329.n22 a_5297_1329.n21 0.223132
R465 a_5297_1329.n23 a_5297_1329.n22 0.223132
R466 a_5297_1329.n24 a_5297_1329.n23 0.223132
R467 a_5297_1329.n26 a_5297_1329.n25 0.153263
R468 a_5297_1329.n14 a_5297_1329.n5 0.139053
R469 a_5297_1329.n16 a_5297_1329.n15 0.124842
R470 a_5297_1329.n30 a_5297_1329.n27 0.114452
R471 a_5297_1329.n13 a_5297_1329.n12 0.110632
R472 a_5297_1329.n15 a_5297_1329.n13 0.108263
R473 a_5297_1329.n16 a_5297_1329.n14 0.0940526
R474 a_5297_1329.n25 a_5297_1329.n5 0.0798421
R475 a_5297_1329.n26 a_5297_1329.n24 0.0656316
R476 a_5297_1329.n31 a_5297_1329.n1 0.0365
R477 a_5297_1329.n29 a_5297_1329.n1 0.0365
R478 a_5297_1329.n28 a_5297_1329.n4 0.0189283
R479 a_5297_1329.n29 a_5297_1329.n28 0.0189283
R480 a_5297_1329.n30 a_5297_1329.n2 0.0130643
R481 a_5297_1329.n2 a_5297_1329.n0 0.0130643
R482 vdd.t5 vdd.t30 1159.16
R483 vdd.t2 vdd.t27 1138.89
R484 vdd.t1 vdd.t29 1132.35
R485 vdd.t3 vdd.n9 888.654
R486 vdd.n2 vdd.t1 522.399
R487 vdd.n10 vdd.t3 522.338
R488 vdd.t30 vdd.n0 522.337
R489 vdd.t29 vdd.n1 517.273
R490 vdd.n1 vdd.t26 517.273
R491 vdd.t27 vdd.n8 517.273
R492 vdd.n8 vdd.t5 517.273
R493 vdd.n9 vdd.t2 513.072
R494 vdd.n4 vdd.t22 304.387
R495 vdd.t22 vdd.t25 208.889
R496 vdd.t25 vdd.t11 208.889
R497 vdd.t11 vdd.t17 208.889
R498 vdd.t17 vdd.t7 208.889
R499 vdd.t7 vdd.t18 208.889
R500 vdd.t18 vdd.t23 208.889
R501 vdd.t23 vdd.t10 208.889
R502 vdd.t10 vdd.t13 208.889
R503 vdd.t13 vdd.t20 208.889
R504 vdd.t20 vdd.t14 208.889
R505 vdd.t14 vdd.t21 208.889
R506 vdd.t21 vdd.t8 208.889
R507 vdd.t8 vdd.t12 208.889
R508 vdd.t12 vdd.t19 208.889
R509 vdd.t19 vdd.t6 208.889
R510 vdd.t6 vdd.t15 208.889
R511 vdd.t15 vdd.t24 208.889
R512 vdd.t24 vdd.t9 208.889
R513 vdd.t9 vdd.t16 208.889
R514 vdd.n6 vdd.t0 9.66464
R515 vdd.n14 vdd.n0 7.11612
R516 vdd.n9 vdd.n5 6.96188
R517 vdd.n2 vdd.n1 6.29206
R518 vdd.n0 vdd.t31 5.262
R519 vdd.n10 vdd.t4 5.26126
R520 vdd.n6 vdd.t28 3.69646
R521 vdd.n4 vdd.n3 3.54271
R522 vdd.n8 vdd.n7 3.13374
R523 vdd.n11 vdd.n10 2.43993
R524 vdd.n13 vdd.n3 2.17281
R525 vdd.n12 vdd.n4 2.08974
R526 vdd.n14 vdd.n13 1.68062
R527 vdd.n7 vdd.n6 1.60498
R528 vdd.n3 vdd.n2 0.698
R529 vdd vdd.n14 0.508779
R530 vdd.n7 vdd.n5 0.337689
R531 vdd.n11 vdd.n5 0.248933
R532 vdd.n13 vdd.n12 0.206214
R533 vdd.n12 vdd.n11 0.0067212
R534 clk.n3 clk.t0 35.7254
R535 clk.n0 clk.t6 35.7221
R536 clk.n5 clk.t5 34.1136
R537 clk.n4 clk.t1 30.1393
R538 clk.n1 clk.t4 30.1393
R539 clk.n2 clk.t2 27.1236
R540 clk.n3 clk.t3 15.823
R541 clk.n0 clk.t7 15.8225
R542 clk.n1 clk.n0 10.6732
R543 clk.n4 clk.n3 10.6727
R544 clk.n6 clk.n2 1.52712
R545 clk clk.n6 0.460065
R546 clk.n6 clk.n5 0.281711
R547 clk.n2 clk.n1 0.111676
R548 clk.n5 clk.n4 0.0995311
R549 nclk.n0 nclk.t7 35.0711
R550 nclk.n3 nclk.t1 28.37
R551 nclk.n1 nclk.t6 25.9811
R552 nclk.n3 nclk.t0 25.2836
R553 nclk.n5 nclk.t4 24.2876
R554 nclk.n2 nclk.t3 24.2876
R555 nclk.n4 nclk.t2 19.9399
R556 nclk.n0 nclk.t5 19.5588
R557 nclk.n2 nclk.n1 7.06888
R558 nclk.n5 nclk.n4 7.0647
R559 nclk.n6 nclk.n5 2.40549
R560 nclk.n6 nclk.n2 1.7803
R561 nclk.n4 nclk.n3 0.699125
R562 nclk nclk.n6 0.594832
R563 nclk.n1 nclk.n0 0.381269
C0 vdd nclk 3.21794f
C1 vin a_8034_n1134# 0.23448f
C2 vin clk 0.14184f
C3 a_8039_2775# nclk 0.68724f
C4 vdd a_8039_2775# 0.86692f
C5 a_8034_n1134# a_5904_n1280# 0.91362f
C6 vin a_5944_2887# 0.05684f
C7 vin vout 15.538f
C8 a_8034_n1134# nclk 0.5632f
C9 vdd a_8034_n1134# 0.5497f
C10 clk a_5904_n1280# 0.82417f
C11 clk nclk 2.7322f
C12 clk vdd 2.16069f
C13 a_5904_n1280# vout 0.00174f
C14 a_5944_2887# nclk 0.12006f
C15 vdd a_5944_2887# 0.3862f
C16 vout nclk 0.17473f
C17 vdd vout 1.94401f
C18 clk a_8039_2775# 0.68185f
C19 a_8039_2775# a_5944_2887# 0.87223f
C20 clk a_8034_n1134# 0.65791f
C21 vin a_5904_n1280# 0.02584f
C22 a_8039_2775# vout 0.00196f
C23 vin nclk 1.46575f
C24 vin vdd 1.55731f
C25 a_8034_n1134# vout 0.00218f
C26 clk a_5944_2887# 0.87934f
C27 clk vout 1.05144f
C28 a_5904_n1280# nclk 0.12185f
C29 vdd a_5904_n1280# 0.23322f
C30 vin a_8039_2775# 0.50886f
C31 a_5944_2887# vout 0.00216f
C32 vout vss 5.0405f
C33 vin vss 3.34778f
C34 nclk vss 6.76557f
C35 clk vss 8.65422f
C36 vdd vss 42.44622f
C37 a_8034_n1134# vss 4.47584f
C38 a_5904_n1280# vss 2.55107f
C39 a_8039_2775# vss 2.74753f
C40 a_5944_2887# vss 1.52239f
C41 nclk.t7 vss 0.02839f
C42 nclk.t5 vss 0.1214f
C43 nclk.n0 vss 0.25404f
C44 nclk.t6 vss 0.13476f
C45 nclk.n1 vss 0.48461f
C46 nclk.t3 vss 0.16661f
C47 nclk.n2 vss 0.58828f
C48 nclk.t2 vss 0.12284f
C49 nclk.t1 vss 0.02302f
C50 nclk.t0 vss 0.12928f
C51 nclk.n3 vss 0.48242f
C52 nclk.n4 vss 0.35941f
C53 nclk.t4 vss 0.16661f
C54 nclk.n5 vss 0.7867f
C55 nclk.n6 vss 1.61769f
C56 clk.t2 vss 0.00995f
C57 clk.t7 vss 0.04631f
C58 clk.t6 vss 0.12799f
C59 clk.n0 vss 0.30308f
C60 clk.t4 vss 0.14359f
C61 clk.n1 vss 0.45504f
C62 clk.n2 vss 0.91656f
C63 clk.t5 vss 0.01691f
C64 clk.t3 vss 0.04631f
C65 clk.t0 vss 0.13424f
C66 clk.n3 vss 0.30815f
C67 clk.t1 vss 0.14359f
C68 clk.n4 vss 0.4463f
C69 clk.n5 vss 0.29462f
C70 clk.n6 vss 1.13327f
C71 vdd.t31 vss 0.0142f
C72 vdd.n0 vss 0.15224f
C73 vdd.t26 vss 0.22942f
C74 vdd.n1 vss 0.42947f
C75 vdd.t29 vss 0.22696f
C76 vdd.t1 vss 0.2285f
C77 vdd.n2 vss 0.22685f
C78 vdd.n3 vss -0.36041f
C79 vdd.t16 vss 0.26651f
C80 vdd.t9 vss 0.12402f
C81 vdd.t24 vss 0.12402f
C82 vdd.t15 vss 0.12402f
C83 vdd.t6 vss 0.12402f
C84 vdd.t19 vss 0.12402f
C85 vdd.t12 vss 0.12402f
C86 vdd.t8 vss 0.12402f
C87 vdd.t21 vss 0.12402f
C88 vdd.t14 vss 0.12402f
C89 vdd.t20 vss 0.12402f
C90 vdd.t13 vss 0.12402f
C91 vdd.t10 vss 0.12402f
C92 vdd.t23 vss 0.12402f
C93 vdd.t18 vss 0.12402f
C94 vdd.t7 vss 0.12402f
C95 vdd.t17 vss 0.12402f
C96 vdd.t11 vss 0.12402f
C97 vdd.t25 vss 0.12402f
C98 vdd.t22 vss 0.15299f
C99 vdd.n4 vss 0.25332f
C100 vdd.n5 vss 0.12916f
C101 vdd.t30 vss 0.16775f
C102 vdd.t5 vss 0.21721f
C103 vdd.t0 vss 0.01245f
C104 vdd.t28 vss 0.02277f
C105 vdd.n6 vss 0.06641f
C106 vdd.n7 vss 0.12516f
C107 vdd.n8 vss 0.4275f
C108 vdd.t27 vss 0.22785f
C109 vdd.t2 vss 0.22676f
C110 vdd.n9 vss 0.1651f
C111 vdd.t3 vss 0.13459f
C112 vdd.t4 vss 0.01423f
C113 vdd.n10 vss 0.12899f
C114 vdd.n11 vss 0.09544f
C115 vdd.n12 vss 0.08296f
C116 vdd.n13 vss 1.41613f
C117 vdd.n14 vss 1.34873f
C118 a_5297_1329.t3 vss 0.06571f
C119 a_5297_1329.n0 vss 0.39189f
C120 a_5297_1329.n1 vss 0.21069f
C121 a_5297_1329.t1 vss 0.0657f
C122 a_5297_1329.t2 vss 0.03559f
C123 a_5297_1329.n3 vss 0.15383f
C124 a_5297_1329.n4 vss 0.17358f
C125 a_5297_1329.n5 vss 0.0225f
C126 a_5297_1329.t13 vss 0.08905f
C127 a_5297_1329.t20 vss 0.08877f
C128 a_5297_1329.n6 vss 0.1212f
C129 a_5297_1329.t5 vss 0.08877f
C130 a_5297_1329.n7 vss 0.06522f
C131 a_5297_1329.t14 vss 0.08877f
C132 a_5297_1329.n8 vss 0.06522f
C133 a_5297_1329.t23 vss 0.08877f
C134 a_5297_1329.n9 vss 0.06522f
C135 a_5297_1329.t10 vss 0.08877f
C136 a_5297_1329.n10 vss 0.06522f
C137 a_5297_1329.t17 vss 0.08877f
C138 a_5297_1329.n11 vss 0.06522f
C139 a_5297_1329.t21 vss 0.08877f
C140 a_5297_1329.n12 vss 0.05775f
C141 a_5297_1329.n13 vss 0.02252f
C142 a_5297_1329.t15 vss 0.08877f
C143 a_5297_1329.n14 vss 0.05108f
C144 a_5297_1329.t8 vss 0.08877f
C145 a_5297_1329.n15 vss 0.05107f
C146 a_5297_1329.n16 vss 0.02251f
C147 a_5297_1329.t7 vss 0.08905f
C148 a_5297_1329.t4 vss 0.08877f
C149 a_5297_1329.n17 vss 0.1212f
C150 a_5297_1329.t18 vss 0.08877f
C151 a_5297_1329.n18 vss 0.06522f
C152 a_5297_1329.t12 vss 0.08877f
C153 a_5297_1329.n19 vss 0.06522f
C154 a_5297_1329.t22 vss 0.08877f
C155 a_5297_1329.n20 vss 0.06522f
C156 a_5297_1329.t11 vss 0.08877f
C157 a_5297_1329.n21 vss 0.06522f
C158 a_5297_1329.t6 vss 0.08877f
C159 a_5297_1329.n22 vss 0.06522f
C160 a_5297_1329.t19 vss 0.08877f
C161 a_5297_1329.n23 vss 0.06522f
C162 a_5297_1329.t16 vss 0.08877f
C163 a_5297_1329.n24 vss 0.0548f
C164 a_5297_1329.t9 vss 0.08877f
C165 a_5297_1329.n25 vss 0.0511f
C166 a_5297_1329.n26 vss 0.02246f
C167 a_5297_1329.n27 vss 0.82798f
C168 a_5297_1329.n29 vss 0.21069f
C169 a_5297_1329.n30 vss 0.89507f
C170 a_5297_1329.n31 vss 0.18815f
C171 a_5297_1329.n32 vss 0.15401f
C172 a_5297_1329.t0 vss 0.03559f
C173 vout.n0 vss 0.11453f
C174 vout.t35 vss 0.27416f
C175 vout.t0 vss 0.22981f
C176 vout.n1 vss 0.71753f
C177 vout.t1 vss 0.04819f
C178 vout.t7 vss 0.04819f
C179 vout.n2 vss 0.1478f
C180 vout.t9 vss 0.04819f
C181 vout.t6 vss 0.04819f
C182 vout.n3 vss 0.1478f
C183 vout.t20 vss 0.06047f
C184 vout.t25 vss 0.06047f
C185 vout.n4 vss 0.18419f
C186 vout.n5 vss 0.33623f
C187 vout.n6 vss 0.11453f
C188 vout.t17 vss 0.04819f
C189 vout.t2 vss 0.04819f
C190 vout.n7 vss 0.1478f
C191 vout.t28 vss 0.06047f
C192 vout.t32 vss 0.06047f
C193 vout.n8 vss 0.18419f
C194 vout.n9 vss 0.11405f
C195 vout.n10 vss 0.11453f
C196 vout.t13 vss 0.04819f
C197 vout.t8 vss 0.04819f
C198 vout.n11 vss 0.1478f
C199 vout.t21 vss 0.06047f
C200 vout.t24 vss 0.06047f
C201 vout.n12 vss 0.18419f
C202 vout.t19 vss 0.04819f
C203 vout.t15 vss 0.04819f
C204 vout.n13 vss 0.1478f
C205 vout.t29 vss 0.06047f
C206 vout.t30 vss 0.06047f
C207 vout.n14 vss 0.18419f
C208 vout.n15 vss 0.33623f
C209 vout.n16 vss 0.11453f
C210 vout.t4 vss 0.04819f
C211 vout.t12 vss 0.04819f
C212 vout.n17 vss 0.1478f
C213 vout.t33 vss 0.06047f
C214 vout.t23 vss 0.06047f
C215 vout.n18 vss 0.18419f
C216 vout.n19 vss 0.11405f
C217 vout.n20 vss 0.11453f
C218 vout.t14 vss 0.04819f
C219 vout.t18 vss 0.04819f
C220 vout.n21 vss 0.1478f
C221 vout.t26 vss 0.06047f
C222 vout.t31 vss 0.06047f
C223 vout.n22 vss 0.18419f
C224 vout.t11 vss 0.04819f
C225 vout.t10 vss 0.04819f
C226 vout.n23 vss 0.1478f
C227 vout.t34 vss 0.06047f
C228 vout.t22 vss 0.06047f
C229 vout.n24 vss 0.18419f
C230 vout.n25 vss 0.33623f
C231 vout.n26 vss 0.20378f
C232 vout.t3 vss 0.04819f
C233 vout.t5 vss 0.04819f
C234 vout.n27 vss 0.1478f
C235 vout.t27 vss 0.27416f
C236 vout.t16 vss 0.22981f
C237 vout.n28 vss 0.7161f
C238 vout.n29 vss 0.01235f
C239 vout.n30 vss 0.18821f
C240 vout.n31 vss 0.10764f
C241 vout.n32 vss 0.0834f
C242 vout.n33 vss 0.11453f
C243 vout.n34 vss 0.11453f
C244 vout.n35 vss 0.08768f
C245 vout.n36 vss 0.10336f
C246 vout.n37 vss 0.33623f
C247 vout.n38 vss 0.06772f
C248 vout.n39 vss 0.11453f
C249 vout.n40 vss 0.11453f
C250 vout.n41 vss 0.11453f
C251 vout.n42 vss 0.06629f
C252 vout.n43 vss 0.33623f
C253 vout.n44 vss 0.10479f
C254 vout.n45 vss 0.08625f
C255 vout.n46 vss 0.11453f
C256 vout.n47 vss 0.11453f
C257 vout.n48 vss 0.08483f
C258 vout.n49 vss 0.10621f
C259 vout.n50 vss 0.33623f
C260 vout.n51 vss 0.06487f
C261 vout.n52 vss 0.11453f
C262 vout.n53 vss 0.11453f
C263 vout.n54 vss 0.11453f
C264 vout.n55 vss 0.06914f
C265 vout.n56 vss 0.33623f
C266 vout.n57 vss 0.10193f
C267 vout.n58 vss 0.0891f
C268 vout.n59 vss 0.11453f
C269 vout.n60 vss 0.11453f
C270 vout.n61 vss 0.08197f
C271 vout.n62 vss 0.10906f
C272 vout.n63 vss 0.18821f
C273 vout.n64 vss 0.00998f
C274 vout.n65 vss 1.03825f
C275 vin.t29 vss 0.03501f
C276 vin.t33 vss 0.03501f
C277 vin.n0 vss 0.11039f
C278 vin.n1 vss 0.24938f
C279 vin.n2 vss 0.56095f
C280 vin.t0 vss 0.0279f
C281 vin.t3 vss 0.0279f
C282 vin.n3 vss 0.09482f
C283 vin.t11 vss 0.0279f
C284 vin.t13 vss 0.0279f
C285 vin.n4 vss 0.08775f
C286 vin.n5 vss 0.42927f
C287 vin.n6 vss 0.14616f
C288 vin.n7 vss 0.17167f
C289 vin.t25 vss 0.03501f
C290 vin.t24 vss 0.03501f
C291 vin.n8 vss 0.1098f
C292 vin.n9 vss 0.13551f
C293 vin.n10 vss 0.10895f
C294 vin.n11 vss 0.18708f
C295 vin.n12 vss 0.09794f
C296 vin.n13 vss 0.56095f
C297 vin.t12 vss 0.0279f
C298 vin.t23 vss 0.0279f
C299 vin.n14 vss 0.08775f
C300 vin.n15 vss 0.09867f
C301 vin.t37 vss 0.03501f
C302 vin.t26 vss 0.03501f
C303 vin.n16 vss 0.1098f
C304 vin.n17 vss 0.13551f
C305 vin.n18 vss 0.18268f
C306 vin.n19 vss 0.11775f
C307 vin.t39 vss 0.03501f
C308 vin.t36 vss 0.03501f
C309 vin.n20 vss 0.1098f
C310 vin.n21 vss 0.13551f
C311 vin.n22 vss 0.16287f
C312 vin.n23 vss 0.56095f
C313 vin.n24 vss 0.12294f
C314 vin.n25 vss 0.13756f
C315 vin.t27 vss 0.03501f
C316 vin.t32 vss 0.03501f
C317 vin.n26 vss 0.1098f
C318 vin.n27 vss 0.13551f
C319 vin.n28 vss 0.14306f
C320 vin.n29 vss 0.15737f
C321 vin.t30 vss 0.03501f
C322 vin.t38 vss 0.03501f
C323 vin.n30 vss 0.1098f
C324 vin.n31 vss 0.13551f
C325 vin.n32 vss 0.12325f
C326 vin.n33 vss 0.56095f
C327 vin.t16 vss 0.0279f
C328 vin.t18 vss 0.0279f
C329 vin.n34 vss 0.08775f
C330 vin.n35 vss 0.09867f
C331 vin.n36 vss 0.14616f
C332 vin.n37 vss 0.17718f
C333 vin.t31 vss 0.03501f
C334 vin.t35 vss 0.03501f
C335 vin.n38 vss 0.1098f
C336 vin.n39 vss 0.13551f
C337 vin.n40 vss 0.10344f
C338 vin.n41 vss 0.18708f
C339 vin.t34 vss 0.03501f
C340 vin.t28 vss 0.03501f
C341 vin.n42 vss 0.10993f
C342 vin.n43 vss 0.19921f
C343 vin.t9 vss 0.0279f
C344 vin.t20 vss 0.0279f
C345 vin.n44 vss 0.09482f
C346 vin.t14 vss 0.0279f
C347 vin.t5 vss 0.0279f
C348 vin.n45 vss 0.08775f
C349 vin.n46 vss 0.40949f
C350 vin.n47 vss 0.08082f
C351 vin.n48 vss 0.80447f
C352 vin.n49 vss 0.56095f
C353 vin.n50 vss 0.56095f
C354 vin.n51 vss 0.08082f
C355 vin.t22 vss 0.0279f
C356 vin.t15 vss 0.0279f
C357 vin.n52 vss 0.08775f
C358 vin.n53 vss 0.09867f
C359 vin.n54 vss 0.13842f
C360 vin.n55 vss 0.09629f
C361 vin.n56 vss 0.56095f
C362 vin.n57 vss 0.56095f
C363 vin.n58 vss 0.56095f
C364 vin.n59 vss 0.11177f
C365 vin.t19 vss 0.0279f
C366 vin.t6 vss 0.0279f
C367 vin.n60 vss 0.08775f
C368 vin.n61 vss 0.09867f
C369 vin.n62 vss 0.10747f
C370 vin.n63 vss 0.12724f
C371 vin.n64 vss 0.56095f
C372 vin.n65 vss 0.56095f
C373 vin.n66 vss 0.09199f
C374 vin.n67 vss 0.14272f
C375 vin.t4 vss 0.0279f
C376 vin.t17 vss 0.0279f
C377 vin.n68 vss 0.08775f
C378 vin.n69 vss 0.09867f
C379 vin.n70 vss 0.07652f
C380 vin.n71 vss 0.56095f
C381 vin.n72 vss 0.56095f
C382 vin.n73 vss 0.56095f
C383 vin.n74 vss 0.08511f
C384 vin.t10 vss 0.0279f
C385 vin.t21 vss 0.0279f
C386 vin.n75 vss 0.08775f
C387 vin.n76 vss 0.09867f
C388 vin.n77 vss 0.13412f
C389 vin.n78 vss 0.10059f
C390 vin.n79 vss 0.33987f
C391 vin.t8 vss 0.03377f
C392 vin.n80 vss 0.02402f
C393 vin.n81 vss 0.07312f
C394 vin.n82 vss 0.01096f
C395 vin.t2 vss 0.04956f
C396 vin.n83 vss 0.05404f
C397 vin.n84 vss 0.01144f
C398 vin.n85 vss 0.0749f
C399 vin.n86 vss 0.43758f
C400 vin.t7 vss 0.03062f
C401 vin.t1 vss 0.04956f
C402 vin.n87 vss 0.12703f
C403 a_5673_n171.n2 vss 0.07314f
C404 a_5673_n171.t2 vss 0.02281f
C405 a_5673_n171.t1 vss 0.01236f
C406 a_5673_n171.n3 vss 0.05347f
C407 a_5673_n171.n4 vss 0.00784f
C408 a_5673_n171.t12 vss 0.03818f
C409 a_5673_n171.t17 vss 0.03809f
C410 a_5673_n171.n5 vss 0.04758f
C411 a_5673_n171.t5 vss 0.03809f
C412 a_5673_n171.n6 vss 0.02544f
C413 a_5673_n171.t8 vss 0.03809f
C414 a_5673_n171.n7 vss 0.02544f
C415 a_5673_n171.t13 vss 0.03809f
C416 a_5673_n171.n8 vss 0.02544f
C417 a_5673_n171.t16 vss 0.03809f
C418 a_5673_n171.n9 vss 0.02272f
C419 a_5673_n171.n10 vss 0.00784f
C420 a_5673_n171.t9 vss 0.03809f
C421 a_5673_n171.n11 vss 0.02029f
C422 a_5673_n171.t6 vss 0.03809f
C423 a_5673_n171.n12 vss 0.02029f
C424 a_5673_n171.n13 vss 0.00784f
C425 a_5673_n171.t4 vss 0.03818f
C426 a_5673_n171.t19 vss 0.03809f
C427 a_5673_n171.n14 vss 0.04758f
C428 a_5673_n171.t14 vss 0.03809f
C429 a_5673_n171.n15 vss 0.02544f
C430 a_5673_n171.t11 vss 0.03809f
C431 a_5673_n171.n16 vss 0.02544f
C432 a_5673_n171.t7 vss 0.03809f
C433 a_5673_n171.n17 vss 0.02544f
C434 a_5673_n171.t18 vss 0.03809f
C435 a_5673_n171.n18 vss 0.02544f
C436 a_5673_n171.t15 vss 0.03809f
C437 a_5673_n171.n19 vss 0.02161f
C438 a_5673_n171.t10 vss 0.03809f
C439 a_5673_n171.n20 vss 0.02029f
C440 a_5673_n171.n21 vss 0.00784f
C441 a_5673_n171.n22 vss 0.26925f
C442 a_5673_n171.n23 vss 0.29043f
C443 a_5673_n171.n24 vss 0.07314f
C444 a_5673_n171.n25 vss 0.06532f
C445 a_5673_n171.n26 vss 0.07178f
C446 a_5673_n171.n27 vss 0.06026f
C447 a_5673_n171.t3 vss 0.01236f
C448 a_5673_n171.n28 vss 0.0534f
C449 a_5673_n171.t0 vss 0.02281f
.ends

