** sch_path: /foss/designs/Mosbious_2025_spiking4all/designs/libs/core_AH_neuron/AH_neuron.sch
.subckt AH_neuron vdd Current_in Vout vss
*.PININFO vdd:B vss:B Current_in:B Vout:B
M5 Vout net1 vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M1 net1 Current_in vdd vdd pfet_03v3 L=0.56u W=0.44u nf=1 m=1
M2 Vout net1 vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M3 net1 Current_in vss vss nfet_03v3 L=0.56u W=0.44u nf=1 m=1
M4 Current_in vgl vss vss nfet_03v3 L=2.4u W=0.22u nf=1 m=1
XC1 Current_in Vout cap_mim_1f0fF c_width=1e-6 c_length=1e-6 m=16
XC2 Vout vgl cap_mim_1f0fF c_width=1e-6 c_length=1e-6 m=1
.ends
