* NGSPICE file created from LIF_comp.ext - technology: gf180mcuD

.subckt pfet$16 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$19 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt switch$2 vdd vss out in cntrl
Xpfet$16_0 m2_n331_n296# cntrl vdd vdd pfet$16
Xpfet$16_1 in m2_n331_n296# out vdd pfet$16
Xnfet$19_0 vss cntrl m2_n331_n296# vss nfet$19
Xnfet$19_1 vss cntrl in out nfet$19
.ends

.subckt pfet$8 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$18 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$2 in1 in2 out cntrl vdd vss
Xpfet$8_0 out cntrl in1 vdd pfet$8
Xpfet$8_1 in2 m2_n850_n472# out vdd pfet$8
Xpfet$8_2 m2_n850_n472# cntrl vdd vdd pfet$8
Xnfet$18_0 vss m2_n850_n472# out in1 nfet$18
Xnfet$18_1 vss cntrl in2 out nfet$18
Xnfet$18_2 vss cntrl m2_n850_n472# vss nfet$18
.ends

.subckt nfet$20 a_n256_n198# a_38_n60# a_n84_0# a_138_0#
X0 a_138_0# a_38_n60# a_n84_0# a_n256_n198# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$17 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$1$5 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$3$2 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt pfet$1$10 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt ota_1stage$2 vss vdd vp vn vout
Xnfet$17_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$17
Xnfet$17_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$17
Xnfet$1$5_0 vss vn vout m2_n516_n58# nfet$1$5
Xnfet$3$2_0 m2_n1824_n806# vss vdd vdd nfet$3$2
Xnfet$1$5_1 vss vp m2_n516_n58# m2_n346_983# nfet$1$5
Xpfet$1$10_0 pfet$1$10_1/w_n352_n286# vout vdd m2_n346_983# pfet$1$10
Xpfet$1$10_1 pfet$1$10_1/w_n352_n286# vdd m2_n346_983# m2_n346_983# pfet$1$10
.ends

.subckt ppolyf_u_resistor$2 a_n376_0# a_160_0# a_n132_0#
X0 a_n132_0# a_160_0# a_n376_0# ppolyf_u r_width=0.8u r_length=0.8u
.ends

.subckt pfet w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$7 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt nfet$5 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$3 a_28_n136# a_n92_0# a_94_0# w_n352_n362#
X0 a_94_0# a_28_n136# a_n92_0# w_n352_n362# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
.ends

.subckt nfet$6 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$4 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_2stages vss vdd vn vp pfet_1/w_n352_n286# vout
Xpfet_0 pfet_1/w_n352_n286# m2_196_146# vdd m2_n346_983# pfet
Xpfet_1 pfet_1/w_n352_n286# vdd m2_n346_983# m2_n346_983# pfet
Xnfet$7_0 vss m2_n516_n58# vss vout nfet$7
Xcap_mim_0 vout m2_196_146# cap_mim
Xnfet$5_0 vss vp m2_196_146# m2_n516_n58# nfet$5
Xnfet$5_1 vss vn m2_n516_n58# m2_n346_983# nfet$5
Xpfet$3_0 m2_196_146# vdd vout pfet_1/w_n352_n286# pfet$3
Xnfet$6_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$6
Xnfet$6_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$6
Xnfet$4_0 m2_n1824_n806# vss vdd vdd nfet$4
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt ppolyf_u_resistor a_n376_0# a_160_0# a_n132_0#
X0 a_n132_0# a_160_0# a_n376_0# ppolyf_u r_width=0.8u r_length=0.8u
.ends

.subckt vdiv vss vspike_up vref vspike_down vres vdd
Xppolyf_u_resistor_18 vdd m1_132_n551# vspike_up ppolyf_u_resistor
Xppolyf_u_resistor_17 vdd m1_56_n1479# m1_n236_n977# ppolyf_u_resistor
Xppolyf_u_resistor_19 vdd m1_132_n551# m1_n236_n977# ppolyf_u_resistor
Xppolyf_u_resistor_0 vdd m1_308_n4993# vss ppolyf_u_resistor
Xppolyf_u_resistor_1 vdd m1_56_n4993# vss ppolyf_u_resistor
Xppolyf_u_resistor_2 vdd m1_308_n4993# m1_600_n4492# ppolyf_u_resistor
Xppolyf_u_resistor_3 vdd m1_56_n4993# m1_n236_n4491# ppolyf_u_resistor
Xppolyf_u_resistor_4 vdd vres m1_n236_n4491# ppolyf_u_resistor
Xppolyf_u_resistor_5 vdd vres m1_600_n4492# ppolyf_u_resistor
Xppolyf_u_resistor_20 vdd m1_132_n49# vspike_up ppolyf_u_resistor
Xppolyf_u_resistor_6 vdd m1_132_n3563# vres ppolyf_u_resistor
Xppolyf_u_resistor_21 vdd m1_132_n49# vdd ppolyf_u_resistor
Xppolyf_u_resistor_10 vdd vref m1_600_n2985# ppolyf_u_resistor
Xppolyf_u_resistor_7 vdd m1_132_n3563# vspike_down ppolyf_u_resistor
Xppolyf_u_resistor_11 vdd vref m1_n236_n2985# ppolyf_u_resistor
Xppolyf_u_resistor_8 vdd vspike_down m1_600_n2985# ppolyf_u_resistor
Xppolyf_u_resistor_12 vdd vref m1_n236_n1981# ppolyf_u_resistor
Xppolyf_u_resistor_9 vdd vspike_down m1_n236_n2985# ppolyf_u_resistor
Xppolyf_u_resistor_13 vdd vref m1_600_n1981# ppolyf_u_resistor
Xppolyf_u_resistor_14 vdd m1_56_n1479# m1_n236_n1981# ppolyf_u_resistor
Xppolyf_u_resistor_15 vdd m1_308_n1479# m1_600_n1981# ppolyf_u_resistor
Xppolyf_u_resistor_16 vdd m1_308_n1479# m1_n236_n977# ppolyf_u_resistor
.ends

.subckt nfet$15 a_n84_n2# a_238_0# a_n256_n272# a_38_n132#
X0 a_238_0# a_38_n132# a_n84_n2# a_n256_n272# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=1u
.ends

.subckt nfet$2$4 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$1$7 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$3$5 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$11 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nand$4 Z A B vdd vss
Xnfet$2$4_0 vss B nfet$3$5_0/a_94_0# vss nfet$2$4
Xpfet$1$7_0 B Z vdd vdd pfet$1$7
Xnfet$3$5_0 A Z nfet$3$5_0/a_94_0# vss nfet$3$5
Xpfet$11_0 A vdd vdd Z pfet$11
.ends

.subckt nfet$11 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$13 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt not$1 vss in out vdd
Xnfet$11_0 vss in out vss nfet$11
Xpfet$13_0 out in vdd vdd pfet$13
.ends

.subckt pfet$7 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$8 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt not vss in vdd
Xpfet$7_0 in in vdd vdd pfet$7
Xnfet$8_0 vss in in vss nfet$8
.ends

.subckt nfet$13 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$15 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt switch$1 vss out in cntrl vdd
Xnfet$13_0 vss cntrl m2_n331_n296# vss nfet$13
Xnfet$13_1 vss cntrl in out nfet$13
Xpfet$15_0 m2_n331_n296# cntrl vdd vdd pfet$15
Xpfet$15_1 in m2_n331_n296# out vdd pfet$15
.ends

.subckt pfet$1$8 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt pfet$2$7 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$10 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$1$3 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nor$2 A B vdd m1_n7_n472# Z vss
Xpfet$1$8_0 m1_n7_n472# vdd Z pfet$1$8_0/a_94_0# pfet$1$8
Xpfet$2$7_0 A pfet$1$8_0/a_94_0# vdd vdd pfet$2$7
Xnfet$10_0 vss A Z vss nfet$10
Xnfet$1$3_0 m1_n7_n472# vss Z vss nfet$1$3
.ends

.subckt nfet$16 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.915p pd=4.22u as=0.915p ps=4.22u w=1.5u l=0.28u
.ends

.subckt pfet$14 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$12 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$1 cntrl out in2 in1 vdd vss
Xpfet$14_0 out cntrl in1 vdd pfet$14
Xpfet$14_1 in2 m2_n850_n472# out vdd pfet$14
Xpfet$14_2 m2_n850_n472# cntrl vdd vdd pfet$14
Xnfet$12_0 vss m2_n850_n472# out in1 nfet$12
Xnfet$12_1 vss cntrl in2 out nfet$12
Xnfet$12_2 vss cntrl m2_n850_n472# vss nfet$12
.ends

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt pfet$1$9 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$1$4 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$14 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$3$6 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_1stage$1 vss vdd vp vn vout
Xpfet$1$9_0 pfet$1$9_1/w_n352_n286# vout vdd m2_n346_983# pfet$1$9
Xpfet$1$9_1 pfet$1$9_1/w_n352_n286# vdd m2_n346_983# m2_n346_983# pfet$1$9
Xnfet$1$4_0 vss vn vout m2_n516_n58# nfet$1$4
Xnfet$1$4_1 vss vp m2_n516_n58# m2_n346_983# nfet$1$4
Xnfet$14_0 vss m2_n1824_n806# m2_n1824_n806# vss nfet$14
Xnfet$14_1 vss m2_n1824_n806# vss m2_n516_n58# nfet$14
Xnfet$3$6_0 m2_n1824_n806# vss vdd vdd nfet$3$6
.ends

.subckt nfet$8$1 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt phaseUpulse reward phi_int phi_2 vspike_up vneg vin vspike ota_1stage$1_0/vdd
+ not$1_0/out vdiv_0/vss not_3/vdd not_3/vss vdiv_0/vref
Xvdiv_0 vdiv_0/vss vspike_up vdiv_0/vref vdiv_0/vspike_down vdiv_0/vres not_3/vss
+ vdiv
Xnfet$15_0 ota_1stage$1_0/vp vneg not_3/vss ota_1stage$1_0/vp nfet$15
Xnand$4_0 nand$4_0/Z vin vneg not_3/vdd not_3/vss nand$4
Xnand$4_1 nand$4_1/Z vneg phi_2 not_3/vdd not_3/vss nand$4
Xnot$1_0 not_3/vss phi_int not$1_0/out not_3/vdd not$1
Xnot_0 not_3/vss vneg not_3/vdd not
Xswitch$1_0 not_3/vss vspike switch$1_0/in vneg not_3/vdd switch$1
Xnot_1 not_3/vss vneg not_3/vdd not
Xnot_2 not_3/vss phi_2 not_3/vdd not
Xnor$2_0 phi_2 nor$2_0/B not_3/vdd vneg phi_int not_3/vss nor$2
Xswitch$1_1 not_3/vss vspike vdiv_0/vref phi_2 not_3/vdd switch$1
Xnfet$16_0 not_3/vss not_3/vss not_3/vss ota_1stage$1_0/vp nfet$16
Xnot_3 not_3/vss phi_2 not_3/vdd not
Xswitch$1_2 not_3/vss vspike switch$1_2/in phi_int not_3/vdd switch$1
Xconmutator$1_0 reward vspike not_3/vdd vspike_up not_3/vdd not_3/vss conmutator$1
Xcap_mim$1_0 vneg nand$4_0/Z cap_mim$1
Xota_1stage$1_0 not_3/vss ota_1stage$1_0/vdd ota_1stage$1_0/vp ota_1stage$1_0/vn switch$1_2/in
+ ota_1stage$1
Xcap_mim$1_1 phi_2 nand$4_1/Z cap_mim$1
Xnfet$8$1_0 not_3/vss ota_1stage$1_0/vn ota_1stage$1_0/vn switch$1_2/in nfet$8$1
Xnfet$8$1_2 not_3/vss vneg vdiv_0/vres not_3/vss nfet$8$1
Xnfet$8$1_1 not_3/vss ota_1stage$1_0/vn vdiv_0/vspike_down vdiv_0/vspike_down nfet$8$1
Xnfet$8$1_3 not_3/vss phi_2 vdiv_0/vres not_3/vss nfet$8$1
.ends

.subckt LIF_comp vout
Xswitch$2_0 switch$2_0/vss switch$2_0/vss switch$2_0/out switch$2_0/in switch$2_0/cntrl
+ switch$2
Xconmutator$2_0 conmutator$2_1/in2 switch$2_0/out vout switch$2_0/cntrl switch$2_0/vss
+ switch$2_0/vss conmutator$2
Xnfet$20_0 switch$2_0/vss ota_1stage$2_0/vn switch$2_0/in switch$2_0/out nfet$20
Xconmutator$2_1 switch$2_0/out conmutator$2_1/in2 conmutator$2_1/out conmutator$2_1/cntrl
+ switch$2_0/vss switch$2_0/vss conmutator$2
Xota_1stage$2_0 switch$2_0/vss switch$2_0/vss ota_1stage$2_0/vp ota_1stage$2_0/vn
+ phaseUpulse_0/vin ota_1stage$2
Xconmutator$2_2 switch$2_0/out switch$2_0/vss ota_1stage$2_0/vp switch$2_0/cntrl switch$2_0/vss
+ switch$2_0/vss conmutator$2
Xppolyf_u_resistor$2_0 switch$2_0/vss ota_1stage$2_0/vn switch$2_0/vss ppolyf_u_resistor$2
Xppolyf_u_resistor$2_1 switch$2_0/vss ota_1stage$2_0/vn m1_2167_4433# ppolyf_u_resistor$2
Xppolyf_u_resistor$2_2 switch$2_0/vss switch$2_0/vss m1_2167_4433# ppolyf_u_resistor$2
Xppolyf_u_resistor$2_3 switch$2_0/vss switch$2_0/vss ppolyf_u_resistor$2_3/a_n132_0#
+ ppolyf_u_resistor$2
Xppolyf_u_resistor$2_4 switch$2_0/vss ota_1stage$2_0/vn switch$2_0/vss ppolyf_u_resistor$2
Xota_2stages_0 switch$2_0/vss switch$2_0/vss switch$2_0/in ota_2stages_0/vp switch$2_0/vss
+ switch$2_0/out ota_2stages
Xcap_mim$3_0 conmutator$2_1/out switch$2_0/in cap_mim$3
XphaseUpulse_0 phaseUpulse_0/reward phaseUpulse_0/phi_int phaseUpulse_0/phi_2 phaseUpulse_0/vspike_up
+ phaseUpulse_0/vneg phaseUpulse_0/vin phaseUpulse_0/vspike switch$2_0/vss switch$2_0/cntrl
+ switch$2_0/vss switch$2_0/vss switch$2_0/vss conmutator$2_1/in2 phaseUpulse
.ends

