* NGSPICE file created from LIF_comp.ext - technology: gf180mcuD

.subckt LIF_comp_pex vdd vss vin v_rew vout
X0 a_n1388_602# ota_1stage$2_0.vout vss.t6 vss.t5 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X1 vspike a_3544_2068# v_ref vdd.t40 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X2 vss.t44 v_rew.t0 a_n872_2246# vss.t43 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X3 vss.t75 phi_fire.t2 a_8075_6021# vss.t74 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X4 v_th phaseUpulse_0.vspike_down phaseUpulse_0.vspike_down vss.t30 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X5 vspike a_2248_2068# phaseUpulse_0.vrefrac vdd.t25 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X6 phaseUpulse_0.vspike_up vdd.t6 vdd.t7 vss.t36 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X7 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.not$1_3.in vdd.t69 vdd.t68 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X8 vdd.t15 vdd.t14 a_6164_1900# vss.t32 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X9 a_2583_6804# v_th ota_1stage$2_0.vout vss.t52 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X10 phaseUpulse_0.phi_2 phaseUpulse_0.monostable_0.not$1_0.in vdd.t44 vdd.t43 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X11 vdd.t42 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.nand$1_0.Z vdd.t41 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X12 vss.t22 phaseUpulse_0.phi_2 a_2248_2068# vss.t21 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X13 vdd.t5 a_2521_8244# ota_1stage$2_0.vout vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X14 a_2328_3444# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp a_2266_4884# vss.t87 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X15 vin.t0 a_8811_n132# vmem.t1 vdd.t32 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X16 vss.t77 phi_fire.t3 a_8827_1078# vss.t76 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X17 vss.t15 phaseUpulse_0.phi_1 a_952_2068# vss.t14 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X18 v_ref a_8827_1078# conmutator$1_2.out vdd.t20 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X19 vdd.t48 v_rew.t1 a_n872_2246# vdd.t47 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X20 phaseUpulse_0.phi_1 phaseUpulse_0.vneg vdd.t3 vdd.t2 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X21 v_ref a_9352_5200# vout.t2 vss.t66 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X22 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vspike_down phaseUpulse_0.vspike_down vss.t29 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X23 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_1 vdd.t31 vdd.t30 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X24 a_7562_3851# a_7562_3851# vdd.t24 vdd.t23 pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X25 vdd.t13 vdd.t12 a_4045_6672# vss.t33 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X26 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.monostable_0.not$1_1.in cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
X27 a_1251_5604# phaseUpulse_0.vspike_up phaseUpulse_0.vspike_up vss.t0 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X28 conmutator$1_2.out phi_fire.t4 vmem.t6 vdd.t32 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X29 vdd.t1 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.nand$1_1.Z vdd.t0 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X30 vmem.t4 v_th vin.t1 vss.t51 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X31 a_4045_6672# a_4045_6672# vss.t71 vss.t69 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X32 a_3790_3312# a_3790_3312# vss.t65 vss.t63 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X33 vss.t17 v_ref v_ref vss.t16 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X34 a_8190_3623# vmem.t2 cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
X35 v_ref phi_fire.t5 conmutator$1_2.out vss.t27 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X36 vdd.t35 phaseUpulse_0.phi_2 a_2248_2068# vdd.t34 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X37 vss.t57 phaseUpulse_0.phi_int a_3544_2068# vss.t56 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X38 a_9352_5200# phi_fire.t6 vdd.t46 vdd.t45 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X39 vin.t3 conmutator$1_2.out cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
X40 vspike phaseUpulse_0.phi_1 phaseUpulse_0.conmutator_0.out vss.t13 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X41 vmem.t3 a_8190_3623# vdd.t54 vdd.t53 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
X42 vdd.t29 phaseUpulse_0.phi_1 a_952_2068# vdd.t28 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X43 phaseUpulse_0.conmutator_0.out v_rew.t2 phaseUpulse_0.vspike_up vdd.t49 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X44 vss.t50 v_th phaseUpulse_0.monostable_0.not$1_3.in vss.t49 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
X45 phaseUpulse_0.monostable_0.nand$1_1.Z ota_1stage$2_0.vout vdd.t17 vdd.t16 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X46 conmutator$1_2.out a_8827_1078# vmem.t0 vss.t8 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X47 vdd.t37 phi_fire.t7 a_8811_n132# vdd.t36 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X48 phaseUpulse_0.phi_int phaseUpulse_0.phi_1 vss.t12 vss.t11 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X49 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.not$1_3.in vss.t84 vss.t83 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X50 vspike phaseUpulse_0.phi_int v_ref vss.t55 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X51 vdd.t52 a_2266_4884# phaseUpulse_0.vrefrac vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X52 vss.t48 v_th phaseUpulse_0.monostable_0.not$1_1.in vss.t47 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
X53 a_7562_3851# vin.t4 a_6854_3116# vss.t23 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X54 ota_1stage$2_0.vp a_8075_6021# vmem.t9 vss.t61 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X55 ota_1stage$2_0.vp phi_fire.t8 vmem.t8 vdd.t38 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X56 vspike phaseUpulse_0.phi_2 phaseUpulse_0.vrefrac vss.t20 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X57 vdd.t59 phaseUpulse_0.phi_int a_3544_2068# vdd.t58 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X58 phaseUpulse_0.phi_1 phaseUpulse_0.vneg vss.t4 vss.t3 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X59 vdd.t4 a_2521_8244# a_2521_8244# vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X60 a_6854_3116# a_6164_1900# vss.t82 vss.t78 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X61 phaseUpulse_0.conmutator_0.out a_n872_2246# phaseUpulse_0.vspike_up vss.t7 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X62 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.monostable_0.not$1_3.in cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
X63 v_ref phi_fire.t9 vout.t0 vdd.t39 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X64 phi_fire.t0 phaseUpulse_0.phi_int vdd.t57 vdd.t56 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X65 a_1078_602# phaseUpulse_0.phi_1 vss.t10 vss.t9 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X66 vdd.t11 vdd.t10 a_3790_3312# vss.t35 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X67 vmem.t11 a_6164_1900# vss.t81 vss.t80 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X68 vdd.t61 phi_fire.t10 a_8827_1078# vdd.t60 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X69 vdd.t22 a_7562_3851# a_8190_3623# vdd.t21 pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X70 phaseUpulse_0.phi_int phaseUpulse_0.phi_2 a_3544_1172# vdd.t33 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X71 a_6854_3116# vspike a_8190_3623# vss.t31 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X72 vdd.t63 phi_fire.t11 a_8075_6021# vdd.t62 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X73 vss.t79 a_6164_1900# a_6164_1900# vss.t78 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X74 vss.t59 phi_fire.t12 a_8811_n132# vss.t58 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X75 vdd.t50 v_rew.t3 phaseUpulse_0.conmutator_0.out vss.t28 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X76 a_2328_3444# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vrefrac vss.t20 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X77 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vss.t86 vss.t85 nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.28u
X78 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in vdd.t67 vdd.t66 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X79 a_3544_1172# phaseUpulse_0.phi_1 vdd.t27 vdd.t26 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X80 vss.t46 v_th v_th vss.t45 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.8u
X81 vout.t1 phi_fire.t13 vmem.t7 vss.t39 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X82 a_2583_6804# ota_1stage$2_0.vp a_2521_8244# vss.t62 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X83 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.vneg phaseUpulse_0.vneg vss.t2 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=3u
X84 v_ref vdd.t8 vdd.t9 vss.t34 nfet_03v3 ad=0.3355p pd=2.32u as=0.3355p ps=2.32u w=0.55u l=0.28u
X85 vin.t2 phi_fire.t14 vmem.t5 vss.t40 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X86 phi_fire.t1 phaseUpulse_0.phi_int vss.t54 vss.t53 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X87 vdd.t19 a_n872_2246# phaseUpulse_0.conmutator_0.out vdd.t18 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X88 vss.t42 phi_fire.t15 ota_1stage$2_0.vp vss.t41 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X89 vss.t60 a_8075_6021# ota_1stage$2_0.vp vdd.t64 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X90 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vneg a_n1388_602# vss.t1 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X91 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.monostable_0.not$1_0.in a_1078_602# vss.t26 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X92 phaseUpulse_0.vrefrac phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.refractory_0.ota_1stage$1_0.vn vss.t67 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X93 vss.t70 a_4045_6672# a_2583_6804# vss.t69 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X94 vdd.t51 a_2266_4884# a_2266_4884# vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X95 vspike a_952_2068# phaseUpulse_0.conmutator_0.out vdd.t55 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X96 vout.t3 a_9352_5200# vmem.t10 vdd.t65 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X97 vss.t64 a_3790_3312# a_2328_3444# vss.t63 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X98 a_9352_5200# phi_fire.t16 vss.t38 vss.t37 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X99 vss.t19 phaseUpulse_0.phi_2 phaseUpulse_0.phi_int vss.t18 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X100 phaseUpulse_0.phi_2 phaseUpulse_0.monostable_0.not$1_0.in vss.t25 vss.t24 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X101 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in vss.t73 vss.t72 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X102 phaseUpulse_0.vspike_down a_1251_5604# a_1251_5604# vss.t68 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
R0 vss.n386 vss.n150 54624.7
R1 vss.n802 vss.n801 12732.4
R2 vss.n386 vss.n321 6691.18
R3 vss.n769 vss.n321 6665.69
R4 vss.n961 vss.n944 6102.12
R5 vss.n202 vss.n150 5709.8
R6 vss.n1180 vss.n1179 4445.99
R7 vss.n274 vss.t34 3683.33
R8 vss.n940 vss.n937 2942.91
R9 vss.n266 vss.n202 2803.92
R10 vss.n1181 vss.n1180 2749.79
R11 vss.n801 vss.t34 2740.2
R12 vss.t53 vss.n832 1853.46
R13 vss.n761 vss.n760 1853.24
R14 vss.n769 vss.n768 1848.04
R15 vss.n1061 vss.n944 1429.64
R16 vss.n1215 vss.n832 1407.47
R17 vss.n803 vss.n802 1363.73
R18 vss.n1021 vss.n943 1314.21
R19 vss.n255 vss.n215 1305.17
R20 vss.n768 vss.n322 1300
R21 vss.n760 vss.n322 1300
R22 vss.n256 vss.n255 1300
R23 vss.n257 vss.n256 1300
R24 vss.n257 vss.n210 1300
R25 vss.n265 vss.n210 1300
R26 vss.n266 vss.n265 1300
R27 vss.t40 vss.t58 1200
R28 vss.n996 vss.n991 910.816
R29 vss.n997 vss.n996 905.739
R30 vss.n998 vss.n997 905.739
R31 vss.n998 vss.n964 905.739
R32 vss.n1019 vss.n964 905.739
R33 vss.n1020 vss.n1019 905.739
R34 vss.n1021 vss.n1020 905.739
R35 vss.n274 vss.n150 892.158
R36 vss.n1180 vss.n942 851.777
R37 vss.t74 vss.t41 799.899
R38 vss.n1179 vss.t58 781.25
R39 vss.n1062 vss.t40 781.25
R40 vss.t18 vss.n1064 740.376
R41 vss.n1158 vss.t26 740.376
R42 vss.n1140 vss.t1 740.376
R43 vss.n1062 vss.n1061 665.625
R44 vss.n1084 vss.n1065 625.567
R45 vss.n1120 vss.n1101 625.567
R46 vss.n939 vss.n938 570.409
R47 vss.n933 vss.t61 487.5
R48 vss.n940 vss.t37 435.103
R49 vss.n1315 vss.n6 432.521
R50 vss.t7 vss.n674 429.632
R51 vss.t41 vss.n933 414.541
R52 vss.t61 vss.n932 414.541
R53 vss.n983 vss.t76 386.286
R54 vss.n1137 vss.t5 378.729
R55 vss vss.t7 376.401
R56 vss.n1064 vss.t53 367.981
R57 vss.n1065 vss.t11 367.981
R58 vss.n1159 vss.t72 367.981
R59 vss.t72 vss.n1158 367.981
R60 vss.n1101 vss.t9 367.981
R61 vss.n1141 vss.t83 367.981
R62 vss.t83 vss.n1140 367.981
R63 vss.n674 vss.t28 365.334
R64 vss.n937 vss.n932 353.19
R65 vss.t11 vss.t18 317.935
R66 vss.t9 vss.t26 317.935
R67 vss.t5 vss.t1 317.935
R68 vss.n1013 vss.n970 290.378
R69 vss.n1411 vss.n127 286.421
R70 vss.n1404 vss.n135 265.962
R71 vss.n522 vss.n515 265.962
R72 vss.n613 vss.n504 265.962
R73 vss.n725 vss.n724 263.036
R74 vss.t66 vss.n941 250.59
R75 vss.n560 vss.n524 248.427
R76 vss.t76 vss.n942 236.606
R77 vss.n723 vss.n422 223.584
R78 vss.n516 vss.n512 216.278
R79 vss.n629 vss.n471 216.278
R80 vss.n1181 vss.t66 213.088
R81 vss.n941 vss.t39 213.088
R82 vss.n613 vss.n498 210.433
R83 vss.n644 vss.n471 210.433
R84 vss.n1160 vss.n1159 195.766
R85 vss.n1142 vss.n1141 195.766
R86 vss.t39 vss.n940 187.517
R87 vss.t27 vss.n974 186.673
R88 vss.n1396 vss.n803 185.589
R89 vss.n1061 vss.n943 177.596
R90 vss.n321 vss.n320 171.47
R91 vss.t80 vss.n974 162.739
R92 vss.t8 vss.n944 154.762
R93 vss.n1168 vss.n1167 150.137
R94 vss.n1160 vss.n1072 150.137
R95 vss.n1150 vss.n1149 150.137
R96 vss.n1142 vss.n1108 150.137
R97 vss.t87 vss.n135 149.056
R98 vss.n551 vss.t87 149.056
R99 vss.t20 vss.n515 149.056
R100 vss.t20 vss.n516 149.056
R101 vss.n620 vss.t85 149.056
R102 vss.t21 vss.n522 146.133
R103 vss.n620 vss.t14 143.21
R104 vss.n698 vss.n697 143.21
R105 vss.n331 vss.n195 142.452
R106 vss.n703 vss.t2 141.75
R107 vss.n652 vss.t13 137.365
R108 vss.n374 vss.n330 134.537
R109 vss.n777 vss.n294 134.537
R110 vss.n749 vss.n393 134.097
R111 vss.n407 vss.n400 134.097
R112 vss.n735 vss.n407 134.097
R113 vss.n725 vss.n409 134.097
R114 vss.n282 vss.t62 131.899
R115 vss.n954 vss.n945 131.125
R116 vss.n1054 vss.n956 131.125
R117 vss.n1232 vss.n921 131.125
R118 vss.n1054 vss.n954 123.919
R119 vss.n644 vss.t14 122.752
R120 vss.t28 vss.n422 122.752
R121 vss.n560 vss.t21 116.906
R122 vss.n1005 vss.n970 113.279
R123 vss.n749 vss.n387 112.731
R124 vss.n791 vss.t62 109.477
R125 vss.n340 vss.n186 109.477
R126 vss.n1198 vss.n930 109.335
R127 vss.n784 vss.n196 104.201
R128 vss.n291 vss.t52 104.201
R129 vss.n983 vss.t27 103.707
R130 vss.n1084 vss.t24 103.034
R131 vss.n1120 vss.t3 103.034
R132 vss.n724 vss.n723 100.832
R133 vss.n1232 vss.n1215 99.4241
R134 vss.n374 vss.n331 98.925
R135 vss.n784 vss.n195 97.606
R136 vss.t37 vss.n939 92.8576
R137 vss.n938 vss.t74 92.8576
R138 vss.n1168 vss.t24 92.7315
R139 vss.n1150 vss.t3 92.7315
R140 vss.n283 vss.n202 85.7351
R141 vss.n449 vss.n447 84.7577
R142 vss.n1275 vss.n869 82.2561
R143 vss.n1308 vss.n857 82.2561
R144 vss.n1482 vss.n6 82.2561
R145 vss.t2 vss.n440 81.835
R146 vss.n681 vss.n432 80.3737
R147 vss.n1411 vss.t55 78.9124
R148 vss.n504 vss.n494 75.9897
R149 vss.n757 vss.n387 75.1535
R150 vss.t0 vss.n393 75.1535
R151 vss.t0 vss.n400 75.1535
R152 vss.n735 vss.t36 75.1535
R153 vss.t36 vss.n409 75.1535
R154 vss.n1167 vss.t47 75.0684
R155 vss.n1149 vss.t49 75.0684
R156 vss.n651 vss.t67 74.5284
R157 vss.n710 vss.t29 74.5284
R158 vss.t31 vss.n945 73.4875
R159 vss.t23 vss.n956 73.4875
R160 vss.t23 vss.n921 73.4875
R161 vss.t85 vss.n494 73.067
R162 vss.n1199 vss.n1198 72.8897
R163 vss.n457 vss.n456 71.6057
R164 vss.n456 vss.n438 70.1444
R165 vss.n164 vss.n163 68.6975
R166 vss.n681 vss.n680 68.6831
R167 vss.n710 vss.n432 68.6831
R168 vss.t45 vss.n340 67.2692
R169 vss.t30 vss.n777 67.2692
R170 vss.n661 vss.t67 67.2217
R171 vss.n698 vss.n440 67.2217
R172 vss.n1013 vss.t8 65.4153
R173 vss.n869 vss.n857 65.0819
R174 vss.n680 vss.n449 64.2991
R175 vss.n670 vss.t43 64.2991
R176 vss.n357 vss.t45 63.3122
R177 vss.n859 vss.n832 58.3025
R178 vss.n1215 vss.n1214 50.7371
R179 vss.n1239 vss.n904 50.6193
R180 vss.t47 vss.n1166 50.0458
R181 vss.t49 vss.n1148 50.0458
R182 vss.t16 vss.n76 49.9628
R183 vss.n1417 vss.t63 49.9628
R184 vss.n512 vss.n498 49.6857
R185 vss.t56 vss.t69 49.473
R186 vss.n1005 vss.t80 49.4605
R187 vss.n724 vss.n420 48.2244
R188 vss.n1247 vss.t78 46.0998
R189 vss.n1275 vss.t78 46.0998
R190 vss.n1061 vss.t31 40.3463
R191 vss.n859 vss.t32 39.7724
R192 vss.n758 vss.t68 37.577
R193 vss.t68 vss.n757 37.577
R194 vss.n778 vss.t30 36.9323
R195 vss.n1199 vss.t51 36.4451
R196 vss.n1214 vss.t51 36.4451
R197 vss.n1463 vss.n73 32.9954
R198 vss.n1482 vss.n7 32.9931
R199 vss.n1247 vss.n904 31.6373
R200 vss.n271 vss.n150 31.3494
R201 vss.t52 vss.n196 30.3374
R202 vss.n778 vss.n291 30.3374
R203 vss.n172 vss.n165 30.0268
R204 vss.n175 vss.n174 30.0268
R205 vss.n728 vss.n727 30.0268
R206 vss.n730 vss.n410 30.0268
R207 vss.n1262 vss.n868 29.7505
R208 vss.n1274 vss.n871 29.7505
R209 vss.n889 vss.n867 29.7505
R210 vss.n1276 vss.n866 29.7505
R211 vss.n1246 vss.n908 29.7505
R212 vss.n115 vss.n97 29.7505
R213 vss.n1435 vss.n99 29.7505
R214 vss.n1412 vss.n120 29.7505
R215 vss.n116 vss.n96 29.7505
R216 vss.n1419 vss.n1418 29.7505
R217 vss.n1462 vss.n77 29.7505
R218 vss.n1465 vss.n71 29.7505
R219 vss.n246 vss.n233 29.7505
R220 vss.n228 vss.n75 29.7505
R221 vss.n225 vss.n223 29.7505
R222 vss.n985 vss.n975 27.1716
R223 vss.n976 vss.n969 27.1716
R224 vss.n937 vss.n930 27.1553
R225 vss.n602 vss.n511 26.8952
R226 vss.n572 vss.n518 26.8952
R227 vss.n672 vss.n451 26.8952
R228 vss.n627 vss.n483 26.8952
R229 vss.n779 vss.n290 26.8952
R230 vss.n318 vss.n292 26.8952
R231 vss.n1476 vss.t35 26.6658
R232 vss.n991 vss.n947 26.2571
R233 vss.n1481 vss.n8 26.2505
R234 vss.n1477 vss.n9 26.2505
R235 vss.n59 vss.n5 26.2505
R236 vss.n1483 vss.n4 26.2505
R237 vss.n1303 vss.n860 26.2505
R238 vss.n1313 vss.n843 26.2505
R239 vss.n1309 vss.n856 26.2505
R240 vss.n1307 vss.n858 26.2505
R241 vss.n1360 vss.n816 26.2505
R242 vss.n1378 vss.n817 26.2505
R243 vss.n827 vss.n814 26.2505
R244 vss.n1381 vss.n1380 26.2505
R245 vss.n645 vss.n465 25.79
R246 vss.n621 vss.n493 25.79
R247 vss.n596 vss.n503 25.79
R248 vss.n615 vss.n495 25.79
R249 vss.n791 vss.n186 25.0614
R250 vss.n1166 vss.n1072 25.0231
R251 vss.n1148 vss.n1108 25.0231
R252 vss.n1012 vss.n1010 24.1237
R253 vss.n1315 vss.n832 23.9541
R254 vss.n1211 vss.n1210 23.9479
R255 vss.n1206 vss.n1205 23.9479
R256 vss.n1189 vss.n929 23.9479
R257 vss.n1197 vss.n931 23.9479
R258 vss.n716 vss.n421 23.9479
R259 vss.n722 vss.n424 23.9479
R260 vss.n695 vss.n433 23.9479
R261 vss.n637 vss.n462 23.9479
R262 vss.n704 vss.n437 23.9479
R263 vss.n804 vss.n93 23.0224
R264 vss.n1177 vss.n1176 22.1935
R265 vss.n1143 vss.n1111 22.0137
R266 vss.n1129 vss.n1112 22.0137
R267 vss.n1122 vss.n1106 22.0137
R268 vss.n1151 vss.n1104 22.0137
R269 vss.n1161 vss.n1075 22.0137
R270 vss.n1093 vss.n1076 22.0137
R271 vss.n1086 vss.n1070 22.0137
R272 vss.n1169 vss.n1068 22.0137
R273 vss.n1438 vss.n1437 21.063
R274 vss.n1417 vss.n114 21.063
R275 vss.n1404 vss.n127 20.4591
R276 vss.n982 vss.n979 20.0599
R277 vss.n272 vss.n92 19.711
R278 vss.n1239 vss.n913 18.5306
R279 vss.n1176 vss 18.2874
R280 vss.n1320 vss.n0 18.0005
R281 vss.n1487 vss.n1486 18.0005
R282 vss.n551 vss.n524 17.5365
R283 vss.n1023 vss.n1022 17.0173
R284 vss.n373 vss.n337 16.8558
R285 vss.n376 vss.n375 16.8558
R286 vss.n405 vss.n402 16.7637
R287 vss.n736 vss.n405 16.7637
R288 vss.n413 vss.n399 16.7637
R289 vss.n413 vss.n408 16.7637
R290 vss.n743 vss.n394 16.6716
R291 vss.n391 vss.n388 16.5794
R292 vss.n157 vss.n94 16.211
R293 vss.n758 vss.n386 16.21
R294 vss.n1438 vss.n93 14.6953
R295 vss.n1437 vss.t69 14.2055
R296 vss.t63 vss.n118 14.2055
R297 vss.n337 vss.n336 14.0926
R298 vss.n301 vss.n296 14.0926
R299 vss.n770 vss.n301 14.0926
R300 vss.n377 vss.n376 14.0926
R301 vss.n384 vss.n383 14.0926
R302 vss.n761 vss.n384 14.0926
R303 vss.n1215 vss.n913 14.0111
R304 vss.n158 vss.n157 13.8163
R305 vss.n276 vss.n187 13.7242
R306 vss.n793 vss.n151 13.7242
R307 vss.n281 vss.n187 13.3558
R308 vss.n794 vss.n793 13.3558
R309 vss.n790 vss.n187 13.3558
R310 vss.n793 vss.n792 13.3558
R311 vss.n747 vss.n394 13.3558
R312 vss.n161 vss.t17 13.2942
R313 vss.n1248 vss.n903 13.2637
R314 vss.n1226 vss.n907 13.2637
R315 vss.n1032 vss.n952 13.2637
R316 vss.n1033 vss.n911 13.2637
R317 vss.n1219 vss.n906 13.2637
R318 vss.n1037 vss.n1029 13.2637
R319 vss.n1031 vss.n903 13.2637
R320 vss.n1029 vss.n1028 13.2637
R321 vss.n952 vss.n948 13.2637
R322 vss.n1395 vss.n1394 13.2637
R323 vss.n545 vss.n514 13.2637
R324 vss.n521 vss.n517 13.2637
R325 vss.n546 vss.n123 13.2637
R326 vss.n550 vss.n521 13.2637
R327 vss.n543 vss.n132 13.2637
R328 vss.n552 vss.n545 13.2637
R329 vss.n1392 vss.n132 13.2637
R330 vss.n1398 vss.n1397 13.2637
R331 vss.n669 vss.n431 13.2637
R332 vss.n485 vss.n478 13.2637
R333 vss.n222 vss.n221 13.2637
R334 vss.n209 vss.n203 13.2637
R335 vss.n787 vss.n786 13.2637
R336 vss.n231 vss.n209 13.2637
R337 vss.n248 vss.n227 13.2637
R338 vss.n783 vss.n197 13.2637
R339 vss.n284 vss.n200 13.2637
R340 vss.n286 vss.n197 13.2637
R341 vss.n786 vss.n785 13.2637
R342 vss.n1439 vss.n92 13.2637
R343 vss.n157 vss.n152 13.2637
R344 vss.n401 vss.n391 13.2637
R345 vss.n411 vss.n405 13.2637
R346 vss.n414 vss.n413 13.2637
R347 vss.n1476 vss.n58 13.1072
R348 vss.n804 vss.n104 11.7563
R349 vss.n181 vss.t46 11.5442
R350 vss vss.n1181 11.0681
R351 vss.n1008 vss.t81 11.0113
R352 vss.n396 vss.n394 10.5926
R353 vss.n1154 vss.n1101 10.59
R354 vss.n1172 vss.n1065 10.59
R355 vss.n675 vss.n674 10.59
R356 vss.n456 vss.n453 10.59
R357 vss.n580 vss.n512 10.59
R358 vss.n541 vss.n127 10.59
R359 vss.n1182 vss.n941 10.59
R360 vss.n1186 vss.n933 10.59
R361 vss.n1187 vss.n932 10.59
R362 vss.n1006 vss.n1005 10.59
R363 vss.n1177 vss.n1062 10.59
R364 vss.n1231 vss.n1216 10.4483
R365 vss.n1403 vss.n136 10.4483
R366 vss.n254 vss.n216 10.4483
R367 vss.n1064 vss.n1063 10.4005
R368 vss.n1166 vss.n1165 10.4005
R369 vss.n1158 vss.n1157 10.4005
R370 vss.n1148 vss.n1147 10.4005
R371 vss.n1140 vss.n1139 10.4005
R372 vss.n539 vss.n524 10.4005
R373 vss.n594 vss.n494 10.4005
R374 vss.n452 vss.n449 10.4005
R375 vss.n805 vss.n804 10.4005
R376 vss.n938 vss.n935 10.4005
R377 vss.n939 vss.n936 10.4005
R378 vss.n973 vss.n942 10.4005
R379 vss.n1179 vss.n1178 10.4005
R380 vss.n699 vss.n445 10.0887
R381 vss.n688 vss.n687 9.85576
R382 vss.n636 vss.n478 9.85576
R383 vss.n691 vss.n442 9.85576
R384 vss.n369 vss.n337 9.85576
R385 vss.n376 vss.n325 9.85576
R386 vss.n767 vss.n301 9.85576
R387 vss.n384 vss.n323 9.85576
R388 vss.n144 vss.t65 9.54445
R389 vss.n250 vss.t71 9.54445
R390 vss.n919 vss.t79 9.54445
R391 vss.n1366 vss.t64 9.54326
R392 vss.n69 vss.t70 9.54326
R393 vss.n1278 vss.t82 9.54326
R394 vss.n1481 vss.n9 9.39524
R395 vss.n1477 vss.n57 9.39524
R396 vss.n1474 vss.n68 9.39524
R397 vss.n1469 vss.n1468 9.39524
R398 vss.n80 vss.n79 9.39524
R399 vss.n1459 vss.n1458 9.39524
R400 vss.n1455 vss.n1454 9.39524
R401 vss.n1451 vss.n1450 9.39524
R402 vss.n1445 vss.n1444 9.39524
R403 vss.n1483 vss.n5 9.39524
R404 vss.n53 vss.n51 9.39524
R405 vss.n51 vss.n50 9.39524
R406 vss.n47 vss.n46 9.39524
R407 vss.n44 vss.n13 9.39524
R408 vss.n40 vss.n38 9.39524
R409 vss.n36 vss.n15 9.39524
R410 vss.n32 vss.n30 9.39524
R411 vss.n28 vss.n17 9.39524
R412 vss.n24 vss.n22 9.39524
R413 vss.n20 vss.n4 9.39524
R414 vss.n1210 vss.n927 9.39524
R415 vss.n1200 vss.n929 9.39524
R416 vss.n1200 vss.n924 9.39524
R417 vss.n1205 vss.n924 9.39524
R418 vss.n1191 vss.n1189 9.39524
R419 vss.n1197 vss.n925 9.39524
R420 vss.n1213 vss.n925 9.39524
R421 vss.n1301 vss.n1300 9.39524
R422 vss.n1297 vss.n1296 9.39524
R423 vss.n1293 vss.n1292 9.39524
R424 vss.n1289 vss.n1288 9.39524
R425 vss.n1317 vss.n831 9.39524
R426 vss.n838 vss.n829 9.39524
R427 vss.n846 vss.n845 9.39524
R428 vss.n850 vss.n849 9.39524
R429 vss.n852 vss.n842 9.39524
R430 vss.n1309 vss.n843 9.39524
R431 vss.n1284 vss.n1282 9.39524
R432 vss.n1282 vss.n1281 9.39524
R433 vss.n882 vss.n880 9.39524
R434 vss.n884 vss.n879 9.39524
R435 vss.n893 vss.n875 9.39524
R436 vss.n1270 vss.n895 9.39524
R437 vss.n1268 vss.n1267 9.39524
R438 vss.n1259 vss.n900 9.39524
R439 vss.n1257 vss.n1256 9.39524
R440 vss.n1253 vss.n856 9.39524
R441 vss.n1307 vss.n860 9.39524
R442 vss.n1133 vss.n1132 9.39524
R443 vss.n1107 vss.n1106 9.39524
R444 vss.n1126 vss.n1107 9.39524
R445 vss.n1126 vss.n1112 9.39524
R446 vss.n1118 vss.n1116 9.39524
R447 vss.n1151 vss.n1105 9.39524
R448 vss.n1144 vss.n1105 9.39524
R449 vss.n1144 vss.n1143 9.39524
R450 vss.n1097 vss.n1096 9.39524
R451 vss.n1071 vss.n1070 9.39524
R452 vss.n1090 vss.n1071 9.39524
R453 vss.n1090 vss.n1076 9.39524
R454 vss.n1082 vss.n1080 9.39524
R455 vss.n1169 vss.n1069 9.39524
R456 vss.n1162 vss.n1069 9.39524
R457 vss.n1162 vss.n1161 9.39524
R458 vss.n1249 vss.n1248 9.39524
R459 vss.n1249 vss.n868 9.39524
R460 vss.n1264 vss.n871 9.39524
R461 vss.n907 vss.n870 9.39524
R462 vss.n1274 vss.n870 9.39524
R463 vss.n1035 vss.n1032 9.39524
R464 vss.n1035 vss.n1033 9.39524
R465 vss.n906 vss.n905 9.39524
R466 vss.n905 vss.n867 9.39524
R467 vss.n887 vss.n866 9.39524
R468 vss.n1246 vss.n865 9.39524
R469 vss.n1276 vss.n865 9.39524
R470 vss.n1037 vss.n1036 9.39524
R471 vss.n1036 vss.n1031 9.39524
R472 vss.n1023 vss.n946 9.39524
R473 vss.n1028 vss.n946 9.39524
R474 vss.n1060 vss.n947 9.39524
R475 vss.n1060 vss.n948 9.39524
R476 vss.n995 vss.n992 9.39524
R477 vss.n995 vss.n990 9.39524
R478 vss.n999 vss.n990 9.39524
R479 vss.n1004 vss.n975 9.39524
R480 vss.n1004 vss.n976 9.39524
R481 vss.n982 vss.n978 9.39524
R482 vss.n1378 vss.n816 9.39524
R483 vss.n1358 vss.n1357 9.39524
R484 vss.n1357 vss.n819 9.39524
R485 vss.n1353 vss.n1351 9.39524
R486 vss.n1349 vss.n821 9.39524
R487 vss.n1345 vss.n1343 9.39524
R488 vss.n1341 vss.n823 9.39524
R489 vss.n1337 vss.n1335 9.39524
R490 vss.n1333 vss.n825 9.39524
R491 vss.n1329 vss.n1327 9.39524
R492 vss.n1325 vss.n827 9.39524
R493 vss.n1380 vss.n814 9.39524
R494 vss.n1374 vss.n817 9.39524
R495 vss.n1372 vss.n1371 9.39524
R496 vss.n1369 vss.n1365 9.39524
R497 vss.n1432 vss.n1431 9.39524
R498 vss.n1429 vss.n105 9.39524
R499 vss.n1425 vss.n1424 9.39524
R500 vss.n1422 vss.n110 9.39524
R501 vss.n1386 vss.n812 9.39524
R502 vss.n119 vss.n115 9.39524
R503 vss.n1395 vss.n119 9.39524
R504 vss.n98 vss.n97 9.39524
R505 vss.n1416 vss.n99 9.39524
R506 vss.n1416 vss.n120 9.39524
R507 vss.n577 vss.n514 9.39524
R508 vss.n577 vss.n511 9.39524
R509 vss.n570 vss.n569 9.39524
R510 vss.n607 vss.n509 9.39524
R511 vss.n605 vss.n604 9.39524
R512 vss.n576 vss.n517 9.39524
R513 vss.n576 vss.n518 9.39524
R514 vss.n549 vss.n546 9.39524
R515 vss.n550 vss.n549 9.39524
R516 vss.n544 vss.n543 9.39524
R517 vss.n552 vss.n544 9.39524
R518 vss.n117 vss.n116 9.39524
R519 vss.n1392 vss.n117 9.39524
R520 vss.n809 vss.n96 9.39524
R521 vss.n1418 vss.n112 9.39524
R522 vss.n1397 vss.n112 9.39524
R523 vss.n718 vss.n424 9.39524
R524 vss.n709 vss.n433 9.39524
R525 vss.n709 vss.n423 9.39524
R526 vss.n722 vss.n423 9.39524
R527 vss.n694 vss.n688 9.39524
R528 vss.n627 vss.n454 9.39524
R529 vss.n662 vss.n454 9.39524
R530 vss.n663 vss.n662 9.39524
R531 vss.n663 vss.n441 9.39524
R532 vss.n446 vss.n441 9.39524
R533 vss.n450 vss.n446 9.39524
R534 vss.n679 vss.n450 9.39524
R535 vss.n679 vss.n451 9.39524
R536 vss.n639 vss.n636 9.39524
R537 vss.n650 vss.n462 9.39524
R538 vss.n650 vss.n436 9.39524
R539 vss.n704 vss.n436 9.39524
R540 vss.n689 vss.n437 9.39524
R541 vss.n645 vss.n466 9.39524
R542 vss.n642 vss.n474 9.39524
R543 vss.n488 vss.n487 9.39524
R544 vss.n596 vss.n492 9.39524
R545 vss.n621 vss.n492 9.39524
R546 vss.n612 vss.n497 9.39524
R547 vss.n612 vss.n505 9.39524
R548 vss.n582 vss.n581 9.39524
R549 vss.n586 vss.n585 9.39524
R550 vss.n590 vss.n589 9.39524
R551 vss.n592 vss.n503 9.39524
R552 vss.n619 vss.n495 9.39524
R553 vss.n619 vss.n465 9.39524
R554 vss.n219 vss.n77 9.39524
R555 vss.n222 vss.n219 9.39524
R556 vss.n1462 vss.n72 9.39524
R557 vss.n232 vss.n71 9.39524
R558 vss.n246 vss.n232 9.39524
R559 vss.n203 vss.n191 9.39524
R560 vss.n787 vss.n191 9.39524
R561 vss.n230 vss.n228 9.39524
R562 vss.n231 vss.n230 9.39524
R563 vss.n1447 vss.n75 9.39524
R564 vss.n226 vss.n225 9.39524
R565 vss.n248 vss.n226 9.39524
R566 vss.n783 vss.n198 9.39524
R567 vss.n779 vss.n198 9.39524
R568 vss.n285 vss.n284 9.39524
R569 vss.n286 vss.n285 9.39524
R570 vss.n785 vss.n193 9.39524
R571 vss.n292 vss.n193 9.39524
R572 vss.n309 vss.n308 9.39524
R573 vss.n313 vss.n312 9.39524
R574 vss.n317 vss.n306 9.39524
R575 vss.n273 vss.n272 9.39524
R576 vss.n165 vss.n91 9.39524
R577 vss.n1439 vss.n91 9.39524
R578 vss.n176 vss.n175 9.39524
R579 vss.n176 vss.n94 9.39524
R580 vss.n155 vss.n154 9.39524
R581 vss.n799 vss.n152 9.39524
R582 vss.n281 vss.n204 9.39524
R583 vss.n369 vss.n368 9.39524
R584 vss.n790 vss.n188 9.39524
R585 vss.n332 vss.n188 9.39524
R586 vss.n373 vss.n332 9.39524
R587 vss.n336 vss.n295 9.39524
R588 vss.n776 vss.n295 9.39524
R589 vss.n776 vss.n296 9.39524
R590 vss.n770 vss.n302 9.39524
R591 vss.n756 vss.n302 9.39524
R592 vss.n756 vss.n388 9.39524
R593 vss.n767 vss.n766 9.39524
R594 vss.n766 vss.n323 9.39524
R595 vss.n792 vss.n184 9.39524
R596 vss.n326 vss.n184 9.39524
R597 vss.n375 vss.n326 9.39524
R598 vss.n378 vss.n377 9.39524
R599 vss.n378 vss.n293 9.39524
R600 vss.n383 vss.n293 9.39524
R601 vss.n761 vss.n759 9.39524
R602 vss.n759 vss.n385 9.39524
R603 vss.n396 vss.n385 9.39524
R604 vss.n750 vss.n392 9.39524
R605 vss.n741 vss.n401 9.39524
R606 vss.n741 vss.n402 9.39524
R607 vss.n736 vss.n406 9.39524
R608 vss.n727 vss.n406 9.39524
R609 vss.n743 vss.n742 9.39524
R610 vss.n742 vss.n399 9.39524
R611 vss.n734 vss.n408 9.39524
R612 vss.n734 vss.n410 9.39524
R613 vss.n1103 vss.t50 9.08339
R614 vss.n1067 vss.t48 9.08339
R615 vss.n1137 vss.t6 9.00997
R616 vss.n1155 vss.t10 9.00997
R617 vss.n1174 vss.t19 9.00997
R618 vss.n1173 vss.t12 9.00997
R619 vss.n633 vss.n467 9.00379
R620 vss.n1178 vss.t59 8.98866
R621 vss.n973 vss.t77 8.98866
R622 vss.n805 vss.t57 8.98866
R623 vss.n594 vss.t15 8.98866
R624 vss.n452 vss.t44 8.98866
R625 vss.n539 vss.t22 8.98866
R626 vss.n936 vss.t75 8.98866
R627 vss.n935 vss.t38 8.98866
R628 vss.n1139 vss.t84 8.98025
R629 vss.n1147 vss.t4 8.98025
R630 vss.n1157 vss.t73 8.98025
R631 vss.n1063 vss.t54 8.98025
R632 vss.n1165 vss.t25 8.98025
R633 vss.n934 vss.t42 8.8205
R634 vss.t43 vss.t29 8.76849
R635 vss vss.t60 8.53506
R636 vss.n154 vss.n92 7.36892
R637 vss.n750 vss.n391 7.36892
R638 vss.n629 vss.n628 7.30715
R639 vss.n652 vss.n651 7.30715
R640 vss.n661 vss.n457 7.30715
R641 vss.n703 vss.n438 7.30715
R642 vss.n479 vss.n468 7.22053
R643 vss.t33 vss.n7 6.77981
R644 vss.n1308 vss.t32 6.32785
R645 vss.n163 vss.t33 6.32785
R646 vss.n697 vss.n447 5.84582
R647 vss.n979 vss.n971 5.40959
R648 vss.n1010 vss.n971 5.40959
R649 vss.n174 vss.n162 5.22638
R650 vss.n1161 vss.n1074 5.2005
R651 vss.n1161 vss.n1160 5.2005
R652 vss.n1163 vss.n1162 5.2005
R653 vss.n1162 vss.n1072 5.2005
R654 vss.n1073 vss.n1069 5.2005
R655 vss.n1167 vss.n1069 5.2005
R656 vss.n1170 vss.n1169 5.2005
R657 vss.n1169 vss.n1168 5.2005
R658 vss.n1068 vss.n1066 5.2005
R659 vss.n1082 vss.n1081 5.2005
R660 vss.n1080 vss.n1079 5.2005
R661 vss.n1087 vss.n1086 5.2005
R662 vss.n1094 vss.n1093 5.2005
R663 vss.n1096 vss.n1095 5.2005
R664 vss.n1098 vss.n1097 5.2005
R665 vss.n1099 vss.n1075 5.2005
R666 vss.n1092 vss.n1076 5.2005
R667 vss.n1160 vss.n1076 5.2005
R668 vss.n1091 vss.n1090 5.2005
R669 vss.n1090 vss.n1072 5.2005
R670 vss.n1089 vss.n1071 5.2005
R671 vss.n1167 vss.n1071 5.2005
R672 vss.n1088 vss.n1070 5.2005
R673 vss.n1168 vss.n1070 5.2005
R674 vss.n1143 vss.n1110 5.2005
R675 vss.n1143 vss.n1142 5.2005
R676 vss.n1145 vss.n1144 5.2005
R677 vss.n1144 vss.n1108 5.2005
R678 vss.n1109 vss.n1105 5.2005
R679 vss.n1149 vss.n1105 5.2005
R680 vss.n1152 vss.n1151 5.2005
R681 vss.n1151 vss.n1150 5.2005
R682 vss.n1104 vss.n1102 5.2005
R683 vss.n1118 vss.n1117 5.2005
R684 vss.n1116 vss.n1115 5.2005
R685 vss.n1123 vss.n1122 5.2005
R686 vss.n1130 vss.n1129 5.2005
R687 vss.n1132 vss.n1131 5.2005
R688 vss.n1134 vss.n1133 5.2005
R689 vss.n1135 vss.n1111 5.2005
R690 vss.n1128 vss.n1112 5.2005
R691 vss.n1142 vss.n1112 5.2005
R692 vss.n1127 vss.n1126 5.2005
R693 vss.n1126 vss.n1108 5.2005
R694 vss.n1125 vss.n1107 5.2005
R695 vss.n1149 vss.n1107 5.2005
R696 vss.n1124 vss.n1106 5.2005
R697 vss.n1150 vss.n1106 5.2005
R698 vss.n302 vss.n300 5.2005
R699 vss.n758 vss.n302 5.2005
R700 vss.n756 vss.n755 5.2005
R701 vss.n757 vss.n756 5.2005
R702 vss.n754 vss.n388 5.2005
R703 vss.n388 vss.n387 5.2005
R704 vss.n411 vss.n403 5.2005
R705 vss.n415 vss.n414 5.2005
R706 vss.n744 vss.n743 5.2005
R707 vss.n743 vss.n393 5.2005
R708 vss.n742 vss.n398 5.2005
R709 vss.n742 vss.t0 5.2005
R710 vss.n416 vss.n399 5.2005
R711 vss.n400 vss.n399 5.2005
R712 vss.n418 vss.n408 5.2005
R713 vss.n735 vss.n408 5.2005
R714 vss.n734 vss.n733 5.2005
R715 vss.t36 vss.n734 5.2005
R716 vss.n732 vss.n410 5.2005
R717 vss.n410 vss.n409 5.2005
R718 vss.n728 vss.n419 5.2005
R719 vss.n731 vss.n730 5.2005
R720 vss.n401 vss.n389 5.2005
R721 vss.n401 vss.n393 5.2005
R722 vss.n741 vss.n740 5.2005
R723 vss.t0 vss.n741 5.2005
R724 vss.n739 vss.n402 5.2005
R725 vss.n402 vss.n400 5.2005
R726 vss.n737 vss.n736 5.2005
R727 vss.n736 vss.n735 5.2005
R728 vss.n406 vss.n404 5.2005
R729 vss.t36 vss.n406 5.2005
R730 vss.n727 vss.n726 5.2005
R731 vss.n727 vss.n409 5.2005
R732 vss.n747 vss.n746 5.2005
R733 vss.n392 vss.n390 5.2005
R734 vss.n751 vss.n750 5.2005
R735 vss.n750 vss.n749 5.2005
R736 vss.n759 vss.n382 5.2005
R737 vss.n759 vss.n758 5.2005
R738 vss.n395 vss.n385 5.2005
R739 vss.n757 vss.n385 5.2005
R740 vss.n397 vss.n396 5.2005
R741 vss.n396 vss.n387 5.2005
R742 vss.n790 vss.n789 5.2005
R743 vss.n791 vss.n790 5.2005
R744 vss.n190 vss.n188 5.2005
R745 vss.n340 vss.n188 5.2005
R746 vss.n362 vss.n332 5.2005
R747 vss.n332 vss.n330 5.2005
R748 vss.n373 vss.n372 5.2005
R749 vss.n374 vss.n373 5.2005
R750 vss.n336 vss.n335 5.2005
R751 vss.n336 vss.n196 5.2005
R752 vss.n333 vss.n295 5.2005
R753 vss.n295 vss.n291 5.2005
R754 vss.n776 vss.n775 5.2005
R755 vss.n777 vss.n776 5.2005
R756 vss.n774 vss.n296 5.2005
R757 vss.n296 vss.n294 5.2005
R758 vss.n795 vss.n794 5.2005
R759 vss.n204 vss.n182 5.2005
R760 vss.n281 vss.n280 5.2005
R761 vss.n282 vss.n281 5.2005
R762 vss.n365 vss.n325 5.2005
R763 vss.n368 vss.n366 5.2005
R764 vss.n370 vss.n369 5.2005
R765 vss.n369 vss.n195 5.2005
R766 vss.n792 vss.n185 5.2005
R767 vss.n792 vss.n791 5.2005
R768 vss.n327 vss.n184 5.2005
R769 vss.n340 vss.n184 5.2005
R770 vss.n328 vss.n326 5.2005
R771 vss.n330 vss.n326 5.2005
R772 vss.n375 vss.n329 5.2005
R773 vss.n375 vss.n374 5.2005
R774 vss.n377 vss.n324 5.2005
R775 vss.n377 vss.n196 5.2005
R776 vss.n379 vss.n378 5.2005
R777 vss.n378 vss.n291 5.2005
R778 vss.n380 vss.n293 5.2005
R779 vss.n777 vss.n293 5.2005
R780 vss.n383 vss.n381 5.2005
R781 vss.n383 vss.n294 5.2005
R782 vss.n318 vss.n298 5.2005
R783 vss.n317 vss.n316 5.2005
R784 vss.n315 vss.n306 5.2005
R785 vss.n314 vss.n313 5.2005
R786 vss.n312 vss.n311 5.2005
R787 vss.n310 vss.n309 5.2005
R788 vss.n308 vss.n307 5.2005
R789 vss.n290 vss.n289 5.2005
R790 vss.n284 vss.n201 5.2005
R791 vss.n284 vss.n283 5.2005
R792 vss.n285 vss.n199 5.2005
R793 vss.n285 vss.t62 5.2005
R794 vss.n287 vss.n286 5.2005
R795 vss.n286 vss.n186 5.2005
R796 vss.n783 vss.n782 5.2005
R797 vss.n784 vss.n783 5.2005
R798 vss.n781 vss.n198 5.2005
R799 vss.t52 vss.n198 5.2005
R800 vss.n780 vss.n779 5.2005
R801 vss.n779 vss.n778 5.2005
R802 vss.n355 vss.n331 5.2005
R803 vss.n331 vss.n192 5.2005
R804 vss.n297 vss.n292 5.2005
R805 vss.n778 vss.n292 5.2005
R806 vss.n334 vss.n193 5.2005
R807 vss.t52 vss.n193 5.2005
R808 vss.n785 vss.n194 5.2005
R809 vss.n785 vss.n784 5.2005
R810 vss.n788 vss.n787 5.2005
R811 vss.n787 vss.n186 5.2005
R812 vss.n191 vss.n189 5.2005
R813 vss.n191 vss.t62 5.2005
R814 vss.n278 vss.n203 5.2005
R815 vss.n283 vss.n203 5.2005
R816 vss.n771 vss.n770 5.2005
R817 vss.n770 vss.n769 5.2005
R818 vss.n764 vss.n323 5.2005
R819 vss.n760 vss.n323 5.2005
R820 vss.n766 vss.n765 5.2005
R821 vss.n766 vss.n322 5.2005
R822 vss.n767 vss.n299 5.2005
R823 vss.n768 vss.n767 5.2005
R824 vss.n762 vss.n761 5.2005
R825 vss.n465 vss.n464 5.2005
R826 vss.n620 vss.n465 5.2005
R827 vss.n619 vss.n618 5.2005
R828 vss.t85 vss.n619 5.2005
R829 vss.n617 vss.n495 5.2005
R830 vss.n504 vss.n495 5.2005
R831 vss.n616 vss.n615 5.2005
R832 vss.n497 vss.n496 5.2005
R833 vss.n612 vss.n611 5.2005
R834 vss.n613 vss.n612 5.2005
R835 vss.n610 vss.n505 5.2005
R836 vss.n581 vss.n506 5.2005
R837 vss.n583 vss.n582 5.2005
R838 vss.n585 vss.n584 5.2005
R839 vss.n587 vss.n586 5.2005
R840 vss.n589 vss.n588 5.2005
R841 vss.n591 vss.n590 5.2005
R842 vss.n593 vss.n592 5.2005
R843 vss.n598 vss.n503 5.2005
R844 vss.n613 vss.n503 5.2005
R845 vss.n493 vss.n490 5.2005
R846 vss.n489 vss.n488 5.2005
R847 vss.n487 vss.n486 5.2005
R848 vss.n480 vss.n479 5.2005
R849 vss.n631 vss.n630 5.2005
R850 vss.n630 vss.n629 5.2005
R851 vss.n654 vss.n653 5.2005
R852 vss.n653 vss.n652 5.2005
R853 vss.n660 vss.n659 5.2005
R854 vss.n661 vss.n660 5.2005
R855 vss.n657 vss.n656 5.2005
R856 vss.n656 vss.n438 5.2005
R857 vss.n702 vss.n701 5.2005
R858 vss.t2 vss.n702 5.2005
R859 vss.n700 vss.n699 5.2005
R860 vss.n699 vss.n698 5.2005
R861 vss.n686 vss.n685 5.2005
R862 vss.n686 vss.n447 5.2005
R863 vss.n684 vss.n448 5.2005
R864 vss.n680 vss.n448 5.2005
R865 vss.n429 vss.n428 5.2005
R866 vss.n432 vss.n429 5.2005
R867 vss.n644 vss.n472 5.2005
R868 vss.n461 vss.n460 5.2005
R869 vss.n628 vss.n461 5.2005
R870 vss.n655 vss.n458 5.2005
R871 vss.n651 vss.n458 5.2005
R872 vss.n658 vss.n459 5.2005
R873 vss.n459 vss.n457 5.2005
R874 vss.n443 vss.n439 5.2005
R875 vss.n703 vss.n439 5.2005
R876 vss.n683 vss.n682 5.2005
R877 vss.n682 vss.n681 5.2005
R878 vss.n712 vss.n711 5.2005
R879 vss.n711 vss.n710 5.2005
R880 vss.n430 vss.n420 5.2005
R881 vss.n723 vss.n421 5.2005
R882 vss.n692 vss.n691 5.2005
R883 vss.n693 vss.n689 5.2005
R884 vss.n437 vss.n434 5.2005
R885 vss.n440 vss.n437 5.2005
R886 vss.n648 vss.n462 5.2005
R887 vss.n628 vss.n462 5.2005
R888 vss.n650 vss.n649 5.2005
R889 vss.n651 vss.n650 5.2005
R890 vss.n436 vss.n435 5.2005
R891 vss.n457 vss.n436 5.2005
R892 vss.n705 vss.n704 5.2005
R893 vss.n704 vss.n703 5.2005
R894 vss.n637 vss.n475 5.2005
R895 vss.n640 vss.n639 5.2005
R896 vss.n636 vss.n635 5.2005
R897 vss.n636 vss.n471 5.2005
R898 vss.n716 vss.n715 5.2005
R899 vss.n719 vss.n718 5.2005
R900 vss.n720 vss.n424 5.2005
R901 vss.n424 vss.n422 5.2005
R902 vss.n707 vss.n433 5.2005
R903 vss.n681 vss.n433 5.2005
R904 vss.n709 vss.n708 5.2005
R905 vss.n710 vss.n709 5.2005
R906 vss.n425 vss.n423 5.2005
R907 vss.n423 vss.n420 5.2005
R908 vss.n722 vss.n721 5.2005
R909 vss.n723 vss.n722 5.2005
R910 vss.n695 vss.n434 5.2005
R911 vss.n694 vss.n693 5.2005
R912 vss.n692 vss.n688 5.2005
R913 vss.n697 vss.n688 5.2005
R914 vss.n634 vss.n633 5.2005
R915 vss.n476 vss.n474 5.2005
R916 vss.n642 vss.n641 5.2005
R917 vss.n466 vss.n463 5.2005
R918 vss.n646 vss.n645 5.2005
R919 vss.n645 vss.n644 5.2005
R920 vss.n644 vss.n467 5.2005
R921 vss.n482 vss.n468 5.2005
R922 vss.n644 vss.n468 5.2005
R923 vss.n486 vss.n485 5.2005
R924 vss.n489 vss.n483 5.2005
R925 vss.n673 vss.n672 5.2005
R926 vss.n669 vss.n427 5.2005
R927 vss.n677 vss.n451 5.2005
R928 vss.n451 vss.n432 5.2005
R929 vss.n679 vss.n678 5.2005
R930 vss.n680 vss.n679 5.2005
R931 vss.n667 vss.n450 5.2005
R932 vss.n450 vss.n447 5.2005
R933 vss.n666 vss.n446 5.2005
R934 vss.n698 vss.n446 5.2005
R935 vss.n665 vss.n441 5.2005
R936 vss.t2 vss.n441 5.2005
R937 vss.n664 vss.n663 5.2005
R938 vss.n663 vss.n438 5.2005
R939 vss.n662 vss.n455 5.2005
R940 vss.n662 vss.n661 5.2005
R941 vss.n625 vss.n454 5.2005
R942 vss.n652 vss.n454 5.2005
R943 vss.n627 vss.n626 5.2005
R944 vss.n629 vss.n627 5.2005
R945 vss.n622 vss.n621 5.2005
R946 vss.n621 vss.n620 5.2005
R947 vss.n492 vss.n491 5.2005
R948 vss.t85 vss.n492 5.2005
R949 vss.n597 vss.n596 5.2005
R950 vss.n596 vss.n504 5.2005
R951 vss.n1393 vss.n143 5.2005
R952 vss.n1395 vss.n149 5.2005
R953 vss.n1396 vss.n1395 5.2005
R954 vss.n1403 vss.n1402 5.2005
R955 vss.n1404 vss.n1403 5.2005
R956 vss.n1397 vss.n149 5.2005
R957 vss.n1397 vss.n1396 5.2005
R958 vss.n1400 vss.n1399 5.2005
R959 vss.n1406 vss.n1405 5.2005
R960 vss.n1405 vss.n1404 5.2005
R961 vss.n1408 vss.n129 5.2005
R962 vss.n1404 vss.n129 5.2005
R963 vss.n130 vss.n128 5.2005
R964 vss.n1404 vss.n128 5.2005
R965 vss.n147 vss.n146 5.2005
R966 vss.n145 vss.n125 5.2005
R967 vss.n1411 vss.n125 5.2005
R968 vss.n1410 vss.n1409 5.2005
R969 vss.n1411 vss.n1410 5.2005
R970 vss.n1407 vss.n126 5.2005
R971 vss.n1411 vss.n126 5.2005
R972 vss.n602 vss.n601 5.2005
R973 vss.n604 vss.n510 5.2005
R974 vss.n605 vss.n508 5.2005
R975 vss.n608 vss.n607 5.2005
R976 vss.n509 vss.n507 5.2005
R977 vss.n569 vss.n567 5.2005
R978 vss.n570 vss.n566 5.2005
R979 vss.n573 vss.n572 5.2005
R980 vss.n547 vss.n546 5.2005
R981 vss.n546 vss.n135 5.2005
R982 vss.n549 vss.n548 5.2005
R983 vss.n549 vss.t87 5.2005
R984 vss.n550 vss.n519 5.2005
R985 vss.n551 vss.n550 5.2005
R986 vss.n565 vss.n517 5.2005
R987 vss.n517 vss.n515 5.2005
R988 vss.n576 vss.n575 5.2005
R989 vss.t20 vss.n576 5.2005
R990 vss.n574 vss.n518 5.2005
R991 vss.n518 vss.n516 5.2005
R992 vss.n562 vss.n522 5.2005
R993 vss.n527 vss.n522 5.2005
R994 vss.n1413 vss.n1412 5.2005
R995 vss.n1412 vss.n1411 5.2005
R996 vss.n140 vss.n139 5.2005
R997 vss.n142 vss.n141 5.2005
R998 vss.n138 vss.n137 5.2005
R999 vss.n579 vss.n511 5.2005
R1000 vss.n516 vss.n511 5.2005
R1001 vss.n578 vss.n577 5.2005
R1002 vss.n577 vss.t20 5.2005
R1003 vss.n514 vss.n513 5.2005
R1004 vss.n515 vss.n514 5.2005
R1005 vss.n553 vss.n552 5.2005
R1006 vss.n552 vss.n551 5.2005
R1007 vss.n544 vss.n540 5.2005
R1008 vss.t87 vss.n544 5.2005
R1009 vss.n543 vss.n542 5.2005
R1010 vss.n543 vss.n135 5.2005
R1011 vss.n1414 vss.n120 5.2005
R1012 vss.n802 vss.n120 5.2005
R1013 vss.n277 vss.n276 5.2005
R1014 vss.n273 vss.n205 5.2005
R1015 vss.n799 vss.n798 5.2005
R1016 vss.n797 vss.n151 5.2005
R1017 vss.n220 vss.n217 5.2005
R1018 vss.n254 vss.n253 5.2005
R1019 vss.n255 vss.n254 5.2005
R1020 vss.n251 vss.n213 5.2005
R1021 vss.n256 vss.n213 5.2005
R1022 vss.n268 vss.n267 5.2005
R1023 vss.n267 vss.n266 5.2005
R1024 vss.n264 vss.n263 5.2005
R1025 vss.n265 vss.n264 5.2005
R1026 vss.n261 vss.n260 5.2005
R1027 vss.n260 vss.n210 5.2005
R1028 vss.n258 vss.n214 5.2005
R1029 vss.n258 vss.n257 5.2005
R1030 vss.n238 vss.n237 5.2005
R1031 vss.n1416 vss.n1415 5.2005
R1032 vss.t63 vss.n1416 5.2005
R1033 vss.n121 vss.n99 5.2005
R1034 vss.n1417 vss.n99 5.2005
R1035 vss.n148 vss.n119 5.2005
R1036 vss.t63 vss.n119 5.2005
R1037 vss.n115 vss.n113 5.2005
R1038 vss.n1417 vss.n115 5.2005
R1039 vss.n148 vss.n112 5.2005
R1040 vss.t63 vss.n112 5.2005
R1041 vss.n1418 vss.n113 5.2005
R1042 vss.n1418 vss.n1417 5.2005
R1043 vss.n272 vss.n270 5.2005
R1044 vss.n272 vss.n271 5.2005
R1045 vss.n1440 vss.n1439 5.2005
R1046 vss.n1439 vss.n1438 5.2005
R1047 vss.n91 vss.n89 5.2005
R1048 vss.t16 vss.n91 5.2005
R1049 vss.n166 vss.n165 5.2005
R1050 vss.n165 vss.n76 5.2005
R1051 vss.n180 vss.n152 5.2005
R1052 vss.n271 vss.n152 5.2005
R1053 vss.n178 vss.n94 5.2005
R1054 vss.n1438 vss.n94 5.2005
R1055 vss.n177 vss.n176 5.2005
R1056 vss.n176 vss.t16 5.2005
R1057 vss.n175 vss.n160 5.2005
R1058 vss.n175 vss.n76 5.2005
R1059 vss.n159 vss.n158 5.2005
R1060 vss.n155 vss.n153 5.2005
R1061 vss.n154 vss.n90 5.2005
R1062 vss.n154 vss.n114 5.2005
R1063 vss.n246 vss.n245 5.2005
R1064 vss.n247 vss.n246 5.2005
R1065 vss.n235 vss.n232 5.2005
R1066 vss.n232 vss.t69 5.2005
R1067 vss.n234 vss.n71 5.2005
R1068 vss.n93 vss.n71 5.2005
R1069 vss.n1466 vss.n1465 5.2005
R1070 vss.n78 vss.n72 5.2005
R1071 vss.n1462 vss.n1461 5.2005
R1072 vss.n1463 vss.n1462 5.2005
R1073 vss.n249 vss.n222 5.2005
R1074 vss.n247 vss.n222 5.2005
R1075 vss.n219 vss.n218 5.2005
R1076 vss.n219 vss.t69 5.2005
R1077 vss.n224 vss.n77 5.2005
R1078 vss.n93 vss.n77 5.2005
R1079 vss.n249 vss.n248 5.2005
R1080 vss.n248 vss.n247 5.2005
R1081 vss.n226 vss.n218 5.2005
R1082 vss.n226 vss.t69 5.2005
R1083 vss.n225 vss.n224 5.2005
R1084 vss.n225 vss.n93 5.2005
R1085 vss.n223 vss.n83 5.2005
R1086 vss.n1448 vss.n1447 5.2005
R1087 vss.n84 vss.n75 5.2005
R1088 vss.n1463 vss.n75 5.2005
R1089 vss.n259 vss.n212 5.2005
R1090 vss.n259 vss.n118 5.2005
R1091 vss.n262 vss.n211 5.2005
R1092 vss.n211 vss.n118 5.2005
R1093 vss.n208 vss.n207 5.2005
R1094 vss.n208 vss.n118 5.2005
R1095 vss.n244 vss.n233 5.2005
R1096 vss.n233 vss.n118 5.2005
R1097 vss.n239 vss.n236 5.2005
R1098 vss.n242 vss.n241 5.2005
R1099 vss.n231 vss.n206 5.2005
R1100 vss.n247 vss.n231 5.2005
R1101 vss.n230 vss.n229 5.2005
R1102 vss.n230 vss.t69 5.2005
R1103 vss.n228 vss.n88 5.2005
R1104 vss.n228 vss.n93 5.2005
R1105 vss.n1392 vss.n1391 5.2005
R1106 vss.n1396 vss.n1392 5.2005
R1107 vss.n1390 vss.n117 5.2005
R1108 vss.t63 vss.n117 5.2005
R1109 vss.n1389 vss.n116 5.2005
R1110 vss.n1417 vss.n116 5.2005
R1111 vss.n1381 vss.n104 5.2005
R1112 vss.n1435 vss.n1434 5.2005
R1113 vss.n101 vss.n98 5.2005
R1114 vss.n106 vss.n97 5.2005
R1115 vss.n1437 vss.n97 5.2005
R1116 vss.n1420 vss.n1419 5.2005
R1117 vss.n810 vss.n809 5.2005
R1118 vss.n807 vss.n96 5.2005
R1119 vss.n1437 vss.n96 5.2005
R1120 vss.n1387 vss.n1386 5.2005
R1121 vss.n812 vss.n811 5.2005
R1122 vss.n111 vss.n110 5.2005
R1123 vss.n1422 vss.n1421 5.2005
R1124 vss.n1424 vss.n109 5.2005
R1125 vss.n1426 vss.n1425 5.2005
R1126 vss.n1427 vss.n105 5.2005
R1127 vss.n1429 vss.n1428 5.2005
R1128 vss.n1431 vss.n103 5.2005
R1129 vss.n1433 vss.n1432 5.2005
R1130 vss.n1365 vss.n100 5.2005
R1131 vss.n1369 vss.n1368 5.2005
R1132 vss.n1371 vss.n1364 5.2005
R1133 vss.n1372 vss.n1363 5.2005
R1134 vss.n1375 vss.n1374 5.2005
R1135 vss.n1376 vss.n817 5.2005
R1136 vss.n817 vss.n104 5.2005
R1137 vss.n986 vss.n985 5.2005
R1138 vss.n978 vss.n977 5.2005
R1139 vss.n982 vss.n981 5.2005
R1140 vss.n983 vss.n982 5.2005
R1141 vss.n1012 vss.n1011 5.2005
R1142 vss.n1013 vss.n1012 5.2005
R1143 vss.n1016 vss.n1015 5.2005
R1144 vss.n969 vss.n967 5.2005
R1145 vss.n1010 vss.n1009 5.2005
R1146 vss.n1010 vss.n970 5.2005
R1147 vss.n972 vss.n971 5.2005
R1148 vss.t80 vss.n971 5.2005
R1149 vss.n980 vss.n979 5.2005
R1150 vss.n979 vss.n974 5.2005
R1151 vss.n987 vss.n975 5.2005
R1152 vss.n975 vss.n974 5.2005
R1153 vss.n1004 vss.n1003 5.2005
R1154 vss.t80 vss.n1004 5.2005
R1155 vss.n1002 vss.n976 5.2005
R1156 vss.n976 vss.n970 5.2005
R1157 vss.n949 vss.n947 5.2005
R1158 vss.n993 vss.n992 5.2005
R1159 vss.n995 vss.n994 5.2005
R1160 vss.n996 vss.n995 5.2005
R1161 vss.n990 vss.n989 5.2005
R1162 vss.n997 vss.n990 5.2005
R1163 vss.n1000 vss.n999 5.2005
R1164 vss.n999 vss.n998 5.2005
R1165 vss.n1022 vss.n963 5.2005
R1166 vss.n1022 vss.n1021 5.2005
R1167 vss.n968 vss.n962 5.2005
R1168 vss.n1020 vss.n962 5.2005
R1169 vss.n1018 vss.n1017 5.2005
R1170 vss.n1019 vss.n1018 5.2005
R1171 vss.n988 vss.n965 5.2005
R1172 vss.n965 vss.n964 5.2005
R1173 vss.n1024 vss.n1023 5.2005
R1174 vss.n1023 vss.n943 5.2005
R1175 vss.n1033 vss.n909 5.2005
R1176 vss.n1033 vss.n921 5.2005
R1177 vss.n1035 vss.n1034 5.2005
R1178 vss.t23 vss.n1035 5.2005
R1179 vss.n1032 vss.n950 5.2005
R1180 vss.n1032 vss.n956 5.2005
R1181 vss.n1058 vss.n948 5.2005
R1182 vss.n948 vss.n945 5.2005
R1183 vss.n1060 vss.n1059 5.2005
R1184 vss.t31 vss.n1060 5.2005
R1185 vss.n1054 vss.n955 5.2005
R1186 vss.n1055 vss.n1054 5.2005
R1187 vss.n1228 vss.n1227 5.2005
R1188 vss.n1231 vss.n1230 5.2005
R1189 vss.n1232 vss.n1231 5.2005
R1190 vss.n1221 vss.n1220 5.2005
R1191 vss.n1218 vss.n1217 5.2005
R1192 vss.n1225 vss.n1224 5.2005
R1193 vss.n918 vss.n916 5.2005
R1194 vss.n1232 vss.n916 5.2005
R1195 vss.n1236 vss.n917 5.2005
R1196 vss.n1232 vss.n917 5.2005
R1197 vss.n1234 vss.n1233 5.2005
R1198 vss.n1233 vss.n1232 5.2005
R1199 vss.n1031 vss.n1030 5.2005
R1200 vss.n1031 vss.n921 5.2005
R1201 vss.n1036 vss.n1027 5.2005
R1202 vss.n1036 vss.t23 5.2005
R1203 vss.n1038 vss.n1037 5.2005
R1204 vss.n1037 vss.n956 5.2005
R1205 vss.n1028 vss.n1026 5.2005
R1206 vss.n1028 vss.n945 5.2005
R1207 vss.n1025 vss.n946 5.2005
R1208 vss.t31 vss.n946 5.2005
R1209 vss.n1277 vss.n1276 5.2005
R1210 vss.n1276 vss.n1275 5.2005
R1211 vss.n865 vss.n864 5.2005
R1212 vss.t78 vss.n865 5.2005
R1213 vss.n1246 vss.n1245 5.2005
R1214 vss.n1247 vss.n1246 5.2005
R1215 vss.n1244 vss.n908 5.2005
R1216 vss.n1239 vss.n908 5.2005
R1217 vss.n1242 vss.n1241 5.2005
R1218 vss.n1262 vss.n1261 5.2005
R1219 vss.n1265 vss.n1264 5.2005
R1220 vss.n897 vss.n871 5.2005
R1221 vss.n871 vss.n869 5.2005
R1222 vss.n1222 vss.n907 5.2005
R1223 vss.n1247 vss.n907 5.2005
R1224 vss.n872 vss.n870 5.2005
R1225 vss.n870 vss.t78 5.2005
R1226 vss.n1274 vss.n1273 5.2005
R1227 vss.n1275 vss.n1274 5.2005
R1228 vss.n1222 vss.n906 5.2005
R1229 vss.n1247 vss.n906 5.2005
R1230 vss.n905 vss.n872 5.2005
R1231 vss.n905 vss.t78 5.2005
R1232 vss.n1273 vss.n867 5.2005
R1233 vss.n1275 vss.n867 5.2005
R1234 vss.n912 vss.n910 5.2005
R1235 vss.n890 vss.n889 5.2005
R1236 vss.n887 vss.n886 5.2005
R1237 vss.n877 vss.n866 5.2005
R1238 vss.n869 vss.n866 5.2005
R1239 vss.n1223 vss.n914 5.2005
R1240 vss.n1239 vss.n914 5.2005
R1241 vss.n1238 vss.n1237 5.2005
R1242 vss.n1239 vss.n1238 5.2005
R1243 vss.n1235 vss.n915 5.2005
R1244 vss.n1239 vss.n915 5.2005
R1245 vss.n1251 vss.n868 5.2005
R1246 vss.n1275 vss.n868 5.2005
R1247 vss.n1250 vss.n1249 5.2005
R1248 vss.n1249 vss.t78 5.2005
R1249 vss.n1248 vss.n902 5.2005
R1250 vss.n1248 vss.n1247 5.2005
R1251 vss.n1305 vss.n860 5.2005
R1252 vss.n860 vss.n859 5.2005
R1253 vss.n1307 vss.n1306 5.2005
R1254 vss.n1308 vss.n1307 5.2005
R1255 vss.n1286 vss.n858 5.2005
R1256 vss.n1285 vss.n1284 5.2005
R1257 vss.n1282 vss.n861 5.2005
R1258 vss.n1282 vss.n857 5.2005
R1259 vss.n1281 vss.n1280 5.2005
R1260 vss.n880 vss.n863 5.2005
R1261 vss.n882 vss.n881 5.2005
R1262 vss.n885 vss.n884 5.2005
R1263 vss.n879 vss.n876 5.2005
R1264 vss.n891 vss.n875 5.2005
R1265 vss.n893 vss.n892 5.2005
R1266 vss.n895 vss.n873 5.2005
R1267 vss.n1271 vss.n1270 5.2005
R1268 vss.n1268 vss.n874 5.2005
R1269 vss.n1267 vss.n1266 5.2005
R1270 vss.n900 vss.n898 5.2005
R1271 vss.n1260 vss.n1259 5.2005
R1272 vss.n1257 vss.n899 5.2005
R1273 vss.n1256 vss.n1255 5.2005
R1274 vss.n1254 vss.n1253 5.2005
R1275 vss.n856 vss.n855 5.2005
R1276 vss.n857 vss.n856 5.2005
R1277 vss.n1313 vss.n1312 5.2005
R1278 vss.n854 vss.n842 5.2005
R1279 vss.n853 vss.n852 5.2005
R1280 vss.n851 vss.n850 5.2005
R1281 vss.n849 vss.n848 5.2005
R1282 vss.n847 vss.n846 5.2005
R1283 vss.n845 vss.n844 5.2005
R1284 vss.n838 vss.n828 5.2005
R1285 vss.n1319 vss.n829 5.2005
R1286 vss.n1318 vss.n1317 5.2005
R1287 vss.n831 vss.n830 5.2005
R1288 vss.n1288 vss.n1287 5.2005
R1289 vss.n1290 vss.n1289 5.2005
R1290 vss.n1292 vss.n1291 5.2005
R1291 vss.n1294 vss.n1293 5.2005
R1292 vss.n1296 vss.n1295 5.2005
R1293 vss.n1298 vss.n1297 5.2005
R1294 vss.n1300 vss.n1299 5.2005
R1295 vss.n1302 vss.n1301 5.2005
R1296 vss.n1304 vss.n1303 5.2005
R1297 vss.n1311 vss.n843 5.2005
R1298 vss.n859 vss.n843 5.2005
R1299 vss.n1310 vss.n1309 5.2005
R1300 vss.n1309 vss.n1308 5.2005
R1301 vss.n1378 vss.n1377 5.2005
R1302 vss.n1379 vss.n1378 5.2005
R1303 vss.n1362 vss.n816 5.2005
R1304 vss.n816 vss.n58 5.2005
R1305 vss.n1361 vss.n1360 5.2005
R1306 vss.n1358 vss.n818 5.2005
R1307 vss.n1357 vss.n1356 5.2005
R1308 vss.n1357 vss.n7 5.2005
R1309 vss.n1355 vss.n819 5.2005
R1310 vss.n1354 vss.n1353 5.2005
R1311 vss.n1351 vss.n820 5.2005
R1312 vss.n1349 vss.n1348 5.2005
R1313 vss.n1347 vss.n821 5.2005
R1314 vss.n1346 vss.n1345 5.2005
R1315 vss.n1343 vss.n822 5.2005
R1316 vss.n1341 vss.n1340 5.2005
R1317 vss.n1339 vss.n823 5.2005
R1318 vss.n1338 vss.n1337 5.2005
R1319 vss.n1335 vss.n824 5.2005
R1320 vss.n1333 vss.n1332 5.2005
R1321 vss.n1331 vss.n825 5.2005
R1322 vss.n1330 vss.n1329 5.2005
R1323 vss.n1327 vss.n826 5.2005
R1324 vss.n1325 vss.n1324 5.2005
R1325 vss.n1323 vss.n827 5.2005
R1326 vss.n827 vss.n7 5.2005
R1327 vss.n1380 vss.n815 5.2005
R1328 vss.n1380 vss.n1379 5.2005
R1329 vss.n1321 vss.n814 5.2005
R1330 vss.n814 vss.n58 5.2005
R1331 vss.n1211 vss.n913 5.2005
R1332 vss.n1207 vss.n1206 5.2005
R1333 vss.n1208 vss.n927 5.2005
R1334 vss.n1210 vss.n1209 5.2005
R1335 vss.n1210 vss.n904 5.2005
R1336 vss.n1205 vss.n1203 5.2005
R1337 vss.n1205 vss.n913 5.2005
R1338 vss.n172 vss.n171 5.2005
R1339 vss.n55 vss.n8 5.2005
R1340 vss.n54 vss.n53 5.2005
R1341 vss.n51 vss.n10 5.2005
R1342 vss.n51 vss.n6 5.2005
R1343 vss.n50 vss.n49 5.2005
R1344 vss.n48 vss.n47 5.2005
R1345 vss.n46 vss.n12 5.2005
R1346 vss.n44 vss.n43 5.2005
R1347 vss.n42 vss.n13 5.2005
R1348 vss.n41 vss.n40 5.2005
R1349 vss.n38 vss.n14 5.2005
R1350 vss.n36 vss.n35 5.2005
R1351 vss.n34 vss.n15 5.2005
R1352 vss.n33 vss.n32 5.2005
R1353 vss.n30 vss.n16 5.2005
R1354 vss.n28 vss.n27 5.2005
R1355 vss.n26 vss.n17 5.2005
R1356 vss.n25 vss.n24 5.2005
R1357 vss.n22 vss.n18 5.2005
R1358 vss.n20 vss.n19 5.2005
R1359 vss.n4 vss.n2 5.2005
R1360 vss.n6 vss.n4 5.2005
R1361 vss.n1476 vss.n59 5.2005
R1362 vss.n1444 vss.n1443 5.2005
R1363 vss.n1446 vss.n1445 5.2005
R1364 vss.n1450 vss.n1449 5.2005
R1365 vss.n1452 vss.n1451 5.2005
R1366 vss.n1454 vss.n1453 5.2005
R1367 vss.n1456 vss.n1455 5.2005
R1368 vss.n1458 vss.n1457 5.2005
R1369 vss.n1460 vss.n1459 5.2005
R1370 vss.n81 vss.n80 5.2005
R1371 vss.n79 vss.n70 5.2005
R1372 vss.n1468 vss.n1467 5.2005
R1373 vss.n1470 vss.n1469 5.2005
R1374 vss.n1472 vss.n68 5.2005
R1375 vss.n1474 vss.n1473 5.2005
R1376 vss.n57 vss.n56 5.2005
R1377 vss.n1478 vss.n1477 5.2005
R1378 vss.n1477 vss.n1476 5.2005
R1379 vss.n5 vss.n3 5.2005
R1380 vss.n163 vss.n5 5.2005
R1381 vss.n1484 vss.n1483 5.2005
R1382 vss.n1483 vss.n1482 5.2005
R1383 vss.n1481 vss.n1480 5.2005
R1384 vss.n1482 vss.n1481 5.2005
R1385 vss.n1479 vss.n9 5.2005
R1386 vss.n163 vss.n9 5.2005
R1387 vss.n1214 vss.n1213 5.2005
R1388 vss.n1195 vss.n925 5.2005
R1389 vss.n1199 vss.n925 5.2005
R1390 vss.n1197 vss.n1196 5.2005
R1391 vss.n1198 vss.n1197 5.2005
R1392 vss.n1193 vss.n931 5.2005
R1393 vss.n1192 vss.n1191 5.2005
R1394 vss.n1189 vss.n1188 5.2005
R1395 vss.n1189 vss.n930 5.2005
R1396 vss.n1202 vss.n924 5.2005
R1397 vss.n1214 vss.n924 5.2005
R1398 vss.n1201 vss.n1200 5.2005
R1399 vss.n1200 vss.n1199 5.2005
R1400 vss.n929 vss.n928 5.2005
R1401 vss.n1198 vss.n929 5.2005
R1402 vss.n1015 vss.n966 5.15839
R1403 vss.n85 vss.n61 4.93742
R1404 vss.n85 vss.n60 4.93742
R1405 vss.n86 vss.n60 4.93742
R1406 vss.n1385 vss.n1384 4.93742
R1407 vss.n1384 vss.n1383 4.93742
R1408 vss.n1383 vss.n1382 4.93742
R1409 vss.n911 vss.n908 4.61478
R1410 vss.n1412 vss.n123 4.61478
R1411 vss.n233 vss.n200 4.61478
R1412 vss.n628 vss.t13 4.38449
R1413 vss.n1012 vss.n966 4.23734
R1414 vss.n1055 vss.n952 4.17792
R1415 vss.n1029 vss.n955 4.17792
R1416 vss.n562 vss.n521 4.04738
R1417 vss.n545 vss.n527 4.04738
R1418 vss.n355 vss.n197 4.04738
R1419 vss.n786 vss.n192 4.04738
R1420 vss.n357 vss.n330 3.95748
R1421 vss.n477 vss.n468 3.938
R1422 vss.n1463 vss.n76 3.91911
R1423 vss.n247 vss.n114 3.91911
R1424 vss.n271 vss.n118 3.91911
R1425 vss.n630 vss.n478 3.66128
R1426 vss.n1233 vss.n903 3.62288
R1427 vss.n1405 vss.n132 3.62288
R1428 vss.n267 vss.n209 3.62288
R1429 vss.n999 vss.n965 3.38837
R1430 vss.n73 vss.t35 3.2919
R1431 vss.n283 vss.n282 2.63849
R1432 vss.n355 vss.n354 2.6005
R1433 vss.n353 vss.n344 2.6005
R1434 vss.n352 vss.n351 2.6005
R1435 vss.n349 vss.n348 2.6005
R1436 vss.n346 vss.n345 2.6005
R1437 vss.n342 vss.n338 2.6005
R1438 vss.n360 vss.n359 2.6005
R1439 vss.n361 vss.n192 2.6005
R1440 vss.n563 vss.n562 2.6005
R1441 vss.n523 vss.n520 2.6005
R1442 vss.n531 vss.n530 2.6005
R1443 vss.n533 vss.n532 2.6005
R1444 vss.n536 vss.n535 2.6005
R1445 vss.n538 vss.n537 2.6005
R1446 vss.n558 vss.n557 2.6005
R1447 vss.n556 vss.n527 2.6005
R1448 vss.n1040 vss.n955 2.6005
R1449 vss.n1043 vss.n1042 2.6005
R1450 vss.n1045 vss.n1044 2.6005
R1451 vss.n1048 vss.n1047 2.6005
R1452 vss.n1050 vss.n1049 2.6005
R1453 vss.n1052 vss.n1051 2.6005
R1454 vss.n959 vss.n951 2.6005
R1455 vss.n1056 vss.n1055 2.6005
R1456 vss.n1018 vss.n965 2.58746
R1457 vss.n1022 vss.n962 2.58746
R1458 vss.n686 vss.n448 2.52347
R1459 vss.n1018 vss.n966 2.51137
R1460 vss.n711 vss.n431 2.49873
R1461 vss.n258 vss.n213 2.497
R1462 vss.n238 vss.n215 2.48287
R1463 vss.n1475 vss.n1474 2.46896
R1464 vss.n1469 vss.n67 2.46896
R1465 vss.n79 vss.n66 2.46896
R1466 vss.n1459 vss.n65 2.46896
R1467 vss.n1455 vss.n64 2.46896
R1468 vss.n1451 vss.n63 2.46896
R1469 vss.n1445 vss.n62 2.46896
R1470 vss.n86 vss.n59 2.46896
R1471 vss.n52 vss.n8 2.46896
R1472 vss.n50 vss.n11 2.46896
R1473 vss.n46 vss.n45 2.46896
R1474 vss.n39 vss.n13 2.46896
R1475 vss.n38 vss.n37 2.46896
R1476 vss.n31 vss.n15 2.46896
R1477 vss.n30 vss.n29 2.46896
R1478 vss.n23 vss.n17 2.46896
R1479 vss.n22 vss.n21 2.46896
R1480 vss.n1206 vss.n1204 2.46896
R1481 vss.n1190 vss.n931 2.46896
R1482 vss.n1212 vss.n1211 2.46896
R1483 vss.n1301 vss.n833 2.46896
R1484 vss.n1297 vss.n834 2.46896
R1485 vss.n1293 vss.n835 2.46896
R1486 vss.n1289 vss.n836 2.46896
R1487 vss.n837 vss.n831 2.46896
R1488 vss.n1316 vss.n829 2.46896
R1489 vss.n845 vss.n839 2.46896
R1490 vss.n849 vss.n840 2.46896
R1491 vss.n852 vss.n841 2.46896
R1492 vss.n1314 vss.n1313 2.46896
R1493 vss.n1283 vss.n858 2.46896
R1494 vss.n1281 vss.n862 2.46896
R1495 vss.n883 vss.n882 2.46896
R1496 vss.n879 vss.n878 2.46896
R1497 vss.n894 vss.n893 2.46896
R1498 vss.n1270 vss.n1269 2.46896
R1499 vss.n1267 vss.n896 2.46896
R1500 vss.n1259 vss.n1258 2.46896
R1501 vss.n1256 vss.n901 2.46896
R1502 vss.n1133 vss.n1113 2.46896
R1503 vss.n1129 vss.n1114 2.46896
R1504 vss.n1119 vss.n1104 2.46896
R1505 vss.n1122 vss.n1121 2.46896
R1506 vss.n1097 vss.n1077 2.46896
R1507 vss.n1093 vss.n1078 2.46896
R1508 vss.n1083 vss.n1068 2.46896
R1509 vss.n1086 vss.n1085 2.46896
R1510 vss.n1083 vss.n1082 2.46896
R1511 vss.n1085 vss.n1080 2.46896
R1512 vss.n1096 vss.n1078 2.46896
R1513 vss.n1077 vss.n1075 2.46896
R1514 vss.n1119 vss.n1118 2.46896
R1515 vss.n1121 vss.n1116 2.46896
R1516 vss.n1132 vss.n1114 2.46896
R1517 vss.n1113 vss.n1111 2.46896
R1518 vss.n1263 vss.n1262 2.46896
R1519 vss.n889 vss.n888 2.46896
R1520 vss.n1015 vss.n1014 2.46896
R1521 vss.n985 vss.n984 2.46896
R1522 vss.n1360 vss.n1359 2.46896
R1523 vss.n1352 vss.n819 2.46896
R1524 vss.n1351 vss.n1350 2.46896
R1525 vss.n1344 vss.n821 2.46896
R1526 vss.n1343 vss.n1342 2.46896
R1527 vss.n1336 vss.n823 2.46896
R1528 vss.n1335 vss.n1334 2.46896
R1529 vss.n1328 vss.n825 2.46896
R1530 vss.n1327 vss.n1326 2.46896
R1531 vss.n1373 vss.n1372 2.46896
R1532 vss.n1370 vss.n1369 2.46896
R1533 vss.n1432 vss.n102 2.46896
R1534 vss.n1430 vss.n1429 2.46896
R1535 vss.n1425 vss.n108 2.46896
R1536 vss.n1423 vss.n1422 2.46896
R1537 vss.n812 vss.n808 2.46896
R1538 vss.n1382 vss.n1381 2.46896
R1539 vss.n1436 vss.n1435 2.46896
R1540 vss.n571 vss.n570 2.46896
R1541 vss.n568 vss.n509 2.46896
R1542 vss.n606 vss.n605 2.46896
R1543 vss.n603 vss.n602 2.46896
R1544 vss.n1419 vss.n95 2.46896
R1545 vss.n717 vss.n716 2.46896
R1546 vss.n696 vss.n695 2.46896
R1547 vss.n672 vss.n671 2.46896
R1548 vss.n485 vss.n484 2.46896
R1549 vss.n638 vss.n637 2.46896
R1550 vss.n691 vss.n690 2.46896
R1551 vss.n643 vss.n642 2.46896
R1552 vss.n633 vss.n473 2.46896
R1553 vss.n487 vss.n469 2.46896
R1554 vss.n493 vss.n470 2.46896
R1555 vss.n615 vss.n614 2.46896
R1556 vss.n505 vss.n499 2.46896
R1557 vss.n582 vss.n500 2.46896
R1558 vss.n586 vss.n501 2.46896
R1559 vss.n590 vss.n502 2.46896
R1560 vss.n1465 vss.n1464 2.46896
R1561 vss.n223 vss.n74 2.46896
R1562 vss.n308 vss.n303 2.46896
R1563 vss.n312 vss.n304 2.46896
R1564 vss.n306 vss.n305 2.46896
R1565 vss.n319 vss.n318 2.46896
R1566 vss.n276 vss.n275 2.46896
R1567 vss.n173 vss.n172 2.46896
R1568 vss.n158 vss.n156 2.46896
R1569 vss.n800 vss.n799 2.46896
R1570 vss.n794 vss.n183 2.46896
R1571 vss.n367 vss.n325 2.46896
R1572 vss.n748 vss.n747 2.46896
R1573 vss.n729 vss.n728 2.46896
R1574 vss.n414 vss.n412 2.46896
R1575 vss.n412 vss.n411 2.46896
R1576 vss.n730 vss.n729 2.46896
R1577 vss.n748 vss.n392 2.46896
R1578 vss.n204 vss.n183 2.46896
R1579 vss.n368 vss.n367 2.46896
R1580 vss.n319 vss.n317 2.46896
R1581 vss.n313 vss.n305 2.46896
R1582 vss.n309 vss.n304 2.46896
R1583 vss.n303 vss.n290 2.46896
R1584 vss.n614 vss.n497 2.46896
R1585 vss.n581 vss.n499 2.46896
R1586 vss.n585 vss.n500 2.46896
R1587 vss.n589 vss.n501 2.46896
R1588 vss.n592 vss.n502 2.46896
R1589 vss.n488 vss.n470 2.46896
R1590 vss.n479 vss.n469 2.46896
R1591 vss.n690 vss.n689 2.46896
R1592 vss.n639 vss.n638 2.46896
R1593 vss.n718 vss.n717 2.46896
R1594 vss.n696 vss.n694 2.46896
R1595 vss.n474 vss.n473 2.46896
R1596 vss.n643 vss.n466 2.46896
R1597 vss.n484 vss.n483 2.46896
R1598 vss.n671 vss.n669 2.46896
R1599 vss.n604 vss.n603 2.46896
R1600 vss.n607 vss.n606 2.46896
R1601 vss.n569 vss.n568 2.46896
R1602 vss.n572 vss.n571 2.46896
R1603 vss.n275 vss.n273 2.46896
R1604 vss.n800 vss.n151 2.46896
R1605 vss.n156 vss.n155 2.46896
R1606 vss.n1464 vss.n72 2.46896
R1607 vss.n1447 vss.n74 2.46896
R1608 vss.n1436 vss.n98 2.46896
R1609 vss.n809 vss.n95 2.46896
R1610 vss.n1386 vss.n1385 2.46896
R1611 vss.n808 vss.n110 2.46896
R1612 vss.n1424 vss.n1423 2.46896
R1613 vss.n108 vss.n105 2.46896
R1614 vss.n1431 vss.n1430 2.46896
R1615 vss.n1365 vss.n102 2.46896
R1616 vss.n1371 vss.n1370 2.46896
R1617 vss.n1374 vss.n1373 2.46896
R1618 vss.n984 vss.n978 2.46896
R1619 vss.n1014 vss.n969 2.46896
R1620 vss.n1264 vss.n1263 2.46896
R1621 vss.n888 vss.n887 2.46896
R1622 vss.n1284 vss.n1283 2.46896
R1623 vss.n880 vss.n862 2.46896
R1624 vss.n884 vss.n883 2.46896
R1625 vss.n878 vss.n875 2.46896
R1626 vss.n895 vss.n894 2.46896
R1627 vss.n1269 vss.n1268 2.46896
R1628 vss.n900 vss.n896 2.46896
R1629 vss.n1258 vss.n1257 2.46896
R1630 vss.n1253 vss.n901 2.46896
R1631 vss.n1314 vss.n842 2.46896
R1632 vss.n850 vss.n841 2.46896
R1633 vss.n846 vss.n840 2.46896
R1634 vss.n839 vss.n838 2.46896
R1635 vss.n1317 vss.n1316 2.46896
R1636 vss.n1288 vss.n837 2.46896
R1637 vss.n1292 vss.n836 2.46896
R1638 vss.n1296 vss.n835 2.46896
R1639 vss.n1300 vss.n834 2.46896
R1640 vss.n1303 vss.n833 2.46896
R1641 vss.n1359 vss.n1358 2.46896
R1642 vss.n1353 vss.n1352 2.46896
R1643 vss.n1350 vss.n1349 2.46896
R1644 vss.n1345 vss.n1344 2.46896
R1645 vss.n1342 vss.n1341 2.46896
R1646 vss.n1337 vss.n1336 2.46896
R1647 vss.n1334 vss.n1333 2.46896
R1648 vss.n1329 vss.n1328 2.46896
R1649 vss.n1326 vss.n1325 2.46896
R1650 vss.n1204 vss.n927 2.46896
R1651 vss.n174 vss.n173 2.46896
R1652 vss.n53 vss.n52 2.46896
R1653 vss.n47 vss.n11 2.46896
R1654 vss.n45 vss.n44 2.46896
R1655 vss.n40 vss.n39 2.46896
R1656 vss.n37 vss.n36 2.46896
R1657 vss.n32 vss.n31 2.46896
R1658 vss.n29 vss.n28 2.46896
R1659 vss.n24 vss.n23 2.46896
R1660 vss.n21 vss.n20 2.46896
R1661 vss.n1444 vss.n61 2.46896
R1662 vss.n1450 vss.n62 2.46896
R1663 vss.n1454 vss.n63 2.46896
R1664 vss.n1458 vss.n64 2.46896
R1665 vss.n80 vss.n65 2.46896
R1666 vss.n1468 vss.n66 2.46896
R1667 vss.n68 vss.n67 2.46896
R1668 vss.n1475 vss.n57 2.46896
R1669 vss.n1213 vss.n1212 2.46896
R1670 vss.n1191 vss.n1190 2.46896
R1671 vss.n653 vss.n461 2.39979
R1672 vss.n660 vss.n458 2.39979
R1673 vss.n656 vss.n459 2.39979
R1674 vss.n702 vss.n439 2.39979
R1675 vss.n1404 vss.n133 2.09769
R1676 vss.n1404 vss.n134 2.09769
R1677 vss.n1411 vss.n124 2.09769
R1678 vss.n240 vss.n118 2.09769
R1679 vss.n1232 vss.n923 2.09769
R1680 vss.n1232 vss.n922 2.09769
R1681 vss.n1240 vss.n1239 2.09769
R1682 vss.n430 vss.n426 2.07536
R1683 vss.n426 vss.n421 2.07536
R1684 vss.n357 vss.n356 2.05118
R1685 vss.n350 vss.n331 2.05118
R1686 vss.n347 vss.n331 2.05118
R1687 vss.n357 vss.n341 2.05118
R1688 vss.n339 vss.n331 2.05118
R1689 vss.n357 vss.n343 2.05118
R1690 vss.n358 vss.n357 2.05118
R1691 vss.n561 vss.n560 2.05118
R1692 vss.n529 vss.n522 2.05118
R1693 vss.n534 vss.n522 2.05118
R1694 vss.n560 vss.n525 2.05118
R1695 vss.n528 vss.n522 2.05118
R1696 vss.n560 vss.n526 2.05118
R1697 vss.n560 vss.n559 2.05118
R1698 vss.n1041 vss.n954 2.03729
R1699 vss.n1054 vss.n957 2.03729
R1700 vss.n1046 vss.n954 2.03729
R1701 vss.n1054 vss.n958 2.03729
R1702 vss.n960 vss.n954 2.03729
R1703 vss.n1054 vss.n1053 2.03729
R1704 vss.n954 vss.n953 2.03729
R1705 vss.n623 vss.t86 1.94108
R1706 vss.n1486 vss.n1 1.86989
R1707 vss.n482 vss.n481 1.76161
R1708 vss.n1224 vss.n914 1.73826
R1709 vss.n1238 vss.n916 1.73826
R1710 vss.n917 vss.n915 1.73826
R1711 vss.n146 vss.n125 1.73826
R1712 vss.n1410 vss.n128 1.73826
R1713 vss.n129 vss.n126 1.73826
R1714 vss.n259 vss.n258 1.73826
R1715 vss.n260 vss.n211 1.73826
R1716 vss.n264 vss.n208 1.73826
R1717 vss.n481 vss.n472 1.67978
R1718 vss.n481 vss.n467 1.67978
R1719 vss.n1487 vss.n0 1.679
R1720 vss.n714 vss.n426 1.56382
R1721 vss.n1396 vss.n150 1.46183
R1722 vss.n803 vss.t55 1.46183
R1723 vss.n670 vss.n420 1.46183
R1724 vss.n702 vss.n442 1.38566
R1725 vss.n1084 vss.n1083 1.36702
R1726 vss.n1085 vss.n1084 1.36702
R1727 vss.n1159 vss.n1078 1.36702
R1728 vss.n1159 vss.n1077 1.36702
R1729 vss.n1120 vss.n1119 1.36702
R1730 vss.n1121 vss.n1120 1.36702
R1731 vss.n1141 vss.n1114 1.36702
R1732 vss.n1141 vss.n1113 1.36702
R1733 vss.n412 vss.n407 1.36702
R1734 vss.n729 vss.n725 1.36702
R1735 vss.n749 vss.n748 1.36702
R1736 vss.n282 vss.n183 1.36702
R1737 vss.n367 vss.n195 1.36702
R1738 vss.n320 vss.n319 1.36702
R1739 vss.n320 vss.n305 1.36702
R1740 vss.n320 vss.n304 1.36702
R1741 vss.n320 vss.n303 1.36702
R1742 vss.n614 vss.n613 1.36702
R1743 vss.n613 vss.n499 1.36702
R1744 vss.n613 vss.n500 1.36702
R1745 vss.n613 vss.n501 1.36702
R1746 vss.n613 vss.n502 1.36702
R1747 vss.n644 vss.n470 1.36702
R1748 vss.n644 vss.n469 1.36702
R1749 vss.n690 vss.n440 1.36702
R1750 vss.n638 vss.n471 1.36702
R1751 vss.n717 vss.n422 1.36702
R1752 vss.n697 vss.n696 1.36702
R1753 vss.n644 vss.n473 1.36702
R1754 vss.n644 vss.n643 1.36702
R1755 vss.n484 vss.n471 1.36702
R1756 vss.n671 vss.n670 1.36702
R1757 vss.n603 vss.n498 1.36702
R1758 vss.n606 vss.n498 1.36702
R1759 vss.n568 vss.n498 1.36702
R1760 vss.n571 vss.n498 1.36702
R1761 vss.n275 vss.n274 1.36702
R1762 vss.n801 vss.n800 1.36702
R1763 vss.n156 vss.n114 1.36702
R1764 vss.n1464 vss.n1463 1.36702
R1765 vss.n1463 vss.n74 1.36702
R1766 vss.n1382 vss.n813 1.36702
R1767 vss.n1383 vss.n104 1.36702
R1768 vss.n1384 vss.n813 1.36702
R1769 vss.n1385 vss.n104 1.36702
R1770 vss.n1437 vss.n1436 1.36702
R1771 vss.n1437 vss.n95 1.36702
R1772 vss.n808 vss.n104 1.36702
R1773 vss.n1423 vss.n104 1.36702
R1774 vss.n108 vss.n104 1.36702
R1775 vss.n1430 vss.n104 1.36702
R1776 vss.n104 vss.n102 1.36702
R1777 vss.n1370 vss.n104 1.36702
R1778 vss.n1373 vss.n104 1.36702
R1779 vss.n984 vss.n983 1.36702
R1780 vss.n1014 vss.n1013 1.36702
R1781 vss.n1263 vss.n869 1.36702
R1782 vss.n888 vss.n869 1.36702
R1783 vss.n1283 vss.n857 1.36702
R1784 vss.n862 vss.n857 1.36702
R1785 vss.n883 vss.n857 1.36702
R1786 vss.n878 vss.n857 1.36702
R1787 vss.n894 vss.n857 1.36702
R1788 vss.n1269 vss.n857 1.36702
R1789 vss.n896 vss.n857 1.36702
R1790 vss.n1258 vss.n857 1.36702
R1791 vss.n901 vss.n857 1.36702
R1792 vss.n1315 vss.n1314 1.36702
R1793 vss.n1315 vss.n841 1.36702
R1794 vss.n1315 vss.n840 1.36702
R1795 vss.n1315 vss.n839 1.36702
R1796 vss.n1316 vss.n1315 1.36702
R1797 vss.n1315 vss.n837 1.36702
R1798 vss.n1315 vss.n836 1.36702
R1799 vss.n1315 vss.n835 1.36702
R1800 vss.n1315 vss.n834 1.36702
R1801 vss.n1315 vss.n833 1.36702
R1802 vss.n1359 vss.n7 1.36702
R1803 vss.n1352 vss.n7 1.36702
R1804 vss.n1350 vss.n7 1.36702
R1805 vss.n1344 vss.n7 1.36702
R1806 vss.n1342 vss.n7 1.36702
R1807 vss.n1336 vss.n7 1.36702
R1808 vss.n1334 vss.n7 1.36702
R1809 vss.n1328 vss.n7 1.36702
R1810 vss.n1326 vss.n7 1.36702
R1811 vss.n1212 vss.n926 1.36702
R1812 vss.n1204 vss.n904 1.36702
R1813 vss.n173 vss.n164 1.36702
R1814 vss.n52 vss.n6 1.36702
R1815 vss.n11 vss.n6 1.36702
R1816 vss.n45 vss.n6 1.36702
R1817 vss.n39 vss.n6 1.36702
R1818 vss.n37 vss.n6 1.36702
R1819 vss.n31 vss.n6 1.36702
R1820 vss.n29 vss.n6 1.36702
R1821 vss.n23 vss.n6 1.36702
R1822 vss.n21 vss.n6 1.36702
R1823 vss.n87 vss.n86 1.36702
R1824 vss.n1476 vss.n60 1.36702
R1825 vss.n87 vss.n85 1.36702
R1826 vss.n1476 vss.n61 1.36702
R1827 vss.n1476 vss.n62 1.36702
R1828 vss.n1476 vss.n63 1.36702
R1829 vss.n1476 vss.n64 1.36702
R1830 vss.n1476 vss.n65 1.36702
R1831 vss.n1476 vss.n66 1.36702
R1832 vss.n1476 vss.n67 1.36702
R1833 vss.n1476 vss.n1475 1.36702
R1834 vss.n1190 vss.n930 1.36702
R1835 vss.n682 vss.n429 1.36092
R1836 vss.n1220 vss.n1219 1.34665
R1837 vss.n1394 vss.n1393 1.34665
R1838 vss.n221 vss.n220 1.34665
R1839 vss.n320 vss.n294 1.31949
R1840 vss.n682 vss.n448 1.16304
R1841 vss.n711 vss.n429 1.16304
R1842 vss.n959 vss.n953 1.12841
R1843 vss.n1053 vss.n1052 1.12841
R1844 vss.n1049 vss.n960 1.12841
R1845 vss.n1047 vss.n958 1.12841
R1846 vss.n1046 vss.n1045 1.12841
R1847 vss.n1042 vss.n957 1.12841
R1848 vss.n1041 vss.n955 1.12841
R1849 vss.n1042 vss.n1041 1.12841
R1850 vss.n1045 vss.n957 1.12841
R1851 vss.n1047 vss.n1046 1.12841
R1852 vss.n1049 vss.n958 1.12841
R1853 vss.n1052 vss.n960 1.12841
R1854 vss.n1053 vss.n959 1.12841
R1855 vss.n1055 vss.n953 1.12841
R1856 vss.n562 vss.n561 1.10063
R1857 vss.n529 vss.n523 1.10063
R1858 vss.n533 vss.n525 1.10063
R1859 vss.n534 vss.n533 1.10063
R1860 vss.n537 vss.n526 1.10063
R1861 vss.n537 vss.n528 1.10063
R1862 vss.n559 vss.n527 1.10063
R1863 vss.n356 vss.n355 1.10063
R1864 vss.n350 vss.n344 1.10063
R1865 vss.n348 vss.n341 1.10063
R1866 vss.n348 vss.n347 1.10063
R1867 vss.n343 vss.n342 1.10063
R1868 vss.n342 vss.n339 1.10063
R1869 vss.n358 vss.n192 1.10063
R1870 vss.n356 vss.n344 1.10063
R1871 vss.n351 vss.n350 1.10063
R1872 vss.n351 vss.n341 1.10063
R1873 vss.n347 vss.n346 1.10063
R1874 vss.n346 vss.n343 1.10063
R1875 vss.n359 vss.n339 1.10063
R1876 vss.n359 vss.n358 1.10063
R1877 vss.n561 vss.n523 1.10063
R1878 vss.n530 vss.n529 1.10063
R1879 vss.n530 vss.n525 1.10063
R1880 vss.n535 vss.n534 1.10063
R1881 vss.n535 vss.n526 1.10063
R1882 vss.n558 vss.n528 1.10063
R1883 vss.n559 vss.n558 1.10063
R1884 vss.n1176 vss.n0 1.0945
R1885 vss.n477 vss.n472 1.02133
R1886 vss.n1379 vss.n73 1.01315
R1887 vss.n1241 vss.n1240 1.00762
R1888 vss.n1220 vss.n922 1.00762
R1889 vss.n1227 vss.n923 1.00762
R1890 vss.n1399 vss.n134 1.00762
R1891 vss.n137 vss.n124 1.00762
R1892 vss.n1393 vss.n133 1.00762
R1893 vss.n241 vss.n240 1.00762
R1894 vss.n146 vss.n134 1.00762
R1895 vss.n140 vss.n124 1.00762
R1896 vss.n141 vss.n133 1.00762
R1897 vss.n240 vss.n239 1.00762
R1898 vss.n1217 vss.n922 1.00762
R1899 vss.n1224 vss.n923 1.00762
R1900 vss.n1240 vss.n912 1.00762
R1901 vss.n687 vss.n445 0.940429
R1902 vss.n478 vss.n477 0.940429
R1903 vss.n445 vss.n442 0.940429
R1904 vss.n1219 vss.n1216 0.93057
R1905 vss.n1226 vss.n1216 0.93057
R1906 vss.n1398 vss.n136 0.93057
R1907 vss.n1394 vss.n136 0.93057
R1908 vss.n227 vss.n216 0.93057
R1909 vss.n221 vss.n216 0.93057
R1910 vss.n1006 vss.n973 0.784993
R1911 vss.n916 vss.n914 0.759241
R1912 vss.n1238 vss.n917 0.759241
R1913 vss.n1233 vss.n915 0.759241
R1914 vss.n128 vss.n125 0.759241
R1915 vss.n1410 vss.n129 0.759241
R1916 vss.n1405 vss.n126 0.759241
R1917 vss.n260 vss.n259 0.759241
R1918 vss.n264 vss.n211 0.759241
R1919 vss.n267 vss.n208 0.759241
R1920 vss.n1138 vss 0.752
R1921 vss.n170 vss.n169 0.6815
R1922 vss.n1178 vss 0.661349
R1923 vss.n1183 vss.n1182 0.603565
R1924 vss.n1241 vss.n911 0.587913
R1925 vss.n137 vss.n123 0.587913
R1926 vss.n241 vss.n200 0.587913
R1927 vss.n1322 vss.n1320 0.552732
R1928 vss.n1217 vss.n912 0.538962
R1929 vss.n141 vss.n140 0.538962
R1930 vss.n239 vss.n238 0.538962
R1931 vss.t16 vss.n104 0.490327
R1932 vss.n247 vss.t56 0.490327
R1933 vss.n169 vss.n168 0.4895
R1934 vss vss.n1177 0.478625
R1935 vss.n1007 vss.n963 0.470735
R1936 vss.n1486 vss.n1485 0.460625
R1937 vss.n164 vss.n58 0.452454
R1938 vss.n1154 vss.n1153 0.450745
R1939 vss.n1172 vss.n1171 0.450745
R1940 vss.n1175 vss.n1174 0.444875
R1941 vss.n1320 vss.n1319 0.434812
R1942 vss.n981 vss.n980 0.426816
R1943 vss.n934 vss 0.396648
R1944 vss.n732 vss.n731 0.386553
R1945 vss.n738 vss 0.38075
R1946 vss.n1414 vss.n1413 0.379017
R1947 vss.n245 vss.n244 0.379017
R1948 vss.n1245 vss.n1244 0.379017
R1949 vss.n162 vss.n161 0.376364
R1950 vss.n987 vss.n986 0.349842
R1951 vss.n574 vss.n573 0.346289
R1952 vss.n780 vss.n289 0.346289
R1953 vss.n993 vss.n949 0.346289
R1954 vss.n676 vss.n675 0.341167
R1955 vss.n1312 vss.n1311 0.338
R1956 vss.n1479 vss.n1478 0.338
R1957 vss.n1480 vss.n55 0.338
R1958 vss.n1377 vss.n1376 0.338
R1959 vss.n1362 vss.n1361 0.338
R1960 vss.n1305 vss.n1304 0.338
R1961 vss.n1306 vss.n1286 0.338
R1962 vss.n1188 vss.n928 0.308395
R1963 vss.n1207 vss.n1203 0.308395
R1964 vss.n1174 vss 0.307625
R1965 vss.n1440 vss.n90 0.302237
R1966 vss.n753 vss 0.302
R1967 vss.n726 vss.n419 0.29236
R1968 vss.n1130 vss.n1128 0.283526
R1969 vss.n1124 vss.n1123 0.283526
R1970 vss.n1094 vss.n1092 0.283526
R1971 vss.n1088 vss.n1087 0.283526
R1972 vss.n171 vss.n167 0.282239
R1973 vss vss.n1136 0.279745
R1974 vss vss.n1100 0.279745
R1975 vss.n617 vss.n616 0.256026
R1976 vss.n1138 vss 0.255875
R1977 vss.n1156 vss 0.255875
R1978 vss vss.n1175 0.255875
R1979 vss.n167 vss.n166 0.231731
R1980 vss.n1310 vss.n855 0.228708
R1981 vss.n417 vss.n416 0.216026
R1982 vss.n418 vss.n417 0.216026
R1983 vss.n179 vss.n178 0.201292
R1984 vss.n745 vss.n744 0.201292
R1985 vss.n598 vss.n597 0.189336
R1986 vss.n646 vss.n464 0.184872
R1987 vss.n721 vss.n720 0.18296
R1988 vss.n1185 vss.n934 0.182778
R1989 vss vss.n1137 0.179375
R1990 vss vss.n1155 0.179375
R1991 vss vss.n1173 0.179375
R1992 vss.n1057 vss.n950 0.171026
R1993 vss.n1243 vss.n909 0.171026
R1994 vss.n547 vss.n122 0.171026
R1995 vss.n564 vss.n519 0.171026
R1996 vss.n565 vss.n564 0.171026
R1997 vss.n782 vss.n288 0.171026
R1998 vss.n243 vss.n201 0.171026
R1999 vss.n288 vss.n287 0.171026
R2000 vss.n738 vss.n403 0.171026
R2001 vss.n417 vss.n415 0.171026
R2002 vss.n1058 vss.n1057 0.171026
R2003 vss.n1002 vss.n1001 0.171026
R2004 vss.n980 vss.n972 0.164429
R2005 vss.n1009 vss.n972 0.164429
R2006 vss.n1367 vss.n1366 0.161799
R2007 vss.n1471 vss.n69 0.161799
R2008 vss.n1279 vss.n1278 0.161799
R2009 vss.n1155 vss.n1154 0.16025
R2010 vss.n1173 vss.n1172 0.16025
R2011 vss.n168 vss.n3 0.1595
R2012 vss.n1187 vss 0.159214
R2013 vss.n1227 vss.n1226 0.147353
R2014 vss.n1399 vss.n1398 0.147353
R2015 vss.n227 vss.n213 0.147353
R2016 vss.n364 vss.n329 0.146252
R2017 vss.n180 vss.n179 0.145456
R2018 vss.n797 vss.n796 0.145456
R2019 vss.n595 vss.n594 0.144974
R2020 vss.n668 vss.n452 0.144974
R2021 vss.n554 vss.n539 0.144974
R2022 vss.n1183 vss.n936 0.144974
R2023 vss.n1184 vss.n935 0.144974
R2024 vss.n806 vss.n805 0.144974
R2025 vss.n1156 vss 0.143375
R2026 vss.n1139 vss.n1138 0.142605
R2027 vss.n1147 vss.n1146 0.142605
R2028 vss.n1157 vss.n1156 0.142605
R2029 vss.n1175 vss.n1063 0.142605
R2030 vss.n1165 vss.n1164 0.142605
R2031 vss.n166 vss.n89 0.141731
R2032 vss.n796 vss.n181 0.140677
R2033 vss.n1209 vss.n926 0.138068
R2034 vss.n715 vss.n714 0.137512
R2035 vss.n1186 vss.n1185 0.134566
R2036 vss.n675 vss 0.134375
R2037 vss.n1182 vss 0.134375
R2038 vss.n601 vss.n600 0.130763
R2039 vss.n773 vss.n298 0.130763
R2040 vss.n179 vss.n159 0.127211
R2041 vss.n371 vss.n370 0.127211
R2042 vss.n365 vss.n364 0.127211
R2043 vss.n772 vss.n299 0.127211
R2044 vss.n764 vss.n763 0.127211
R2045 vss.n746 vss.n745 0.127211
R2046 vss.n280 vss.n279 0.127211
R2047 vss.n796 vss.n795 0.127211
R2048 vss.n1136 vss.n1135 0.126026
R2049 vss.n1153 vss.n1102 0.126026
R2050 vss.n1100 vss.n1099 0.126026
R2051 vss.n1171 vss.n1066 0.126026
R2052 vss.n630 vss.n461 0.124175
R2053 vss.n653 vss.n458 0.124175
R2054 vss.n660 vss.n459 0.124175
R2055 vss.n656 vss.n439 0.124175
R2056 vss.n1485 vss.n2 0.122474
R2057 vss.n1323 vss.n1322 0.122474
R2058 vss.n364 vss.n324 0.122358
R2059 vss.n763 vss.n381 0.122358
R2060 vss.n763 vss.n762 0.122358
R2061 vss.n745 vss.n397 0.122358
R2062 vss.n752 vss.n389 0.121833
R2063 vss.n739 vss.n738 0.121833
R2064 vss.n738 vss.n737 0.121833
R2065 vss.n1135 vss.n1134 0.121289
R2066 vss.n1134 vss.n1131 0.121289
R2067 vss.n1131 vss.n1130 0.121289
R2068 vss.n1125 vss.n1124 0.121289
R2069 vss.n1127 vss.n1125 0.121289
R2070 vss.n1128 vss.n1127 0.121289
R2071 vss.n1117 vss.n1102 0.121289
R2072 vss.n1117 vss.n1115 0.121289
R2073 vss.n1123 vss.n1115 0.121289
R2074 vss.n1099 vss.n1098 0.121289
R2075 vss.n1098 vss.n1095 0.121289
R2076 vss.n1095 vss.n1094 0.121289
R2077 vss.n1089 vss.n1088 0.121289
R2078 vss.n1091 vss.n1089 0.121289
R2079 vss.n1092 vss.n1091 0.121289
R2080 vss.n1081 vss.n1066 0.121289
R2081 vss.n1081 vss.n1079 0.121289
R2082 vss.n1087 vss.n1079 0.121289
R2083 vss.n1034 vss.n950 0.121289
R2084 vss.n1034 vss.n909 0.121289
R2085 vss.n1311 vss.n1310 0.121289
R2086 vss.n844 vss.n828 0.121289
R2087 vss.n847 vss.n844 0.121289
R2088 vss.n848 vss.n847 0.121289
R2089 vss.n851 vss.n848 0.121289
R2090 vss.n853 vss.n851 0.121289
R2091 vss.n854 vss.n853 0.121289
R2092 vss.n1312 vss.n854 0.121289
R2093 vss.n720 vss.n719 0.121289
R2094 vss.n719 vss.n715 0.121289
R2095 vss.n618 vss.n617 0.121289
R2096 vss.n618 vss.n464 0.121289
R2097 vss.n548 vss.n547 0.121289
R2098 vss.n548 vss.n519 0.121289
R2099 vss.n575 vss.n565 0.121289
R2100 vss.n575 vss.n574 0.121289
R2101 vss.n573 vss.n566 0.121289
R2102 vss.n567 vss.n566 0.121289
R2103 vss.n567 vss.n507 0.121289
R2104 vss.n608 vss.n508 0.121289
R2105 vss.n510 vss.n508 0.121289
R2106 vss.n601 vss.n510 0.121289
R2107 vss.n1193 vss.n1192 0.121289
R2108 vss.n1192 vss.n1188 0.121289
R2109 vss.n1201 vss.n928 0.121289
R2110 vss.n1202 vss.n1201 0.121289
R2111 vss.n1203 vss.n1202 0.121289
R2112 vss.n1209 vss.n1208 0.121289
R2113 vss.n1208 vss.n1207 0.121289
R2114 vss.n307 vss.n289 0.121289
R2115 vss.n310 vss.n307 0.121289
R2116 vss.n311 vss.n310 0.121289
R2117 vss.n314 vss.n311 0.121289
R2118 vss.n315 vss.n314 0.121289
R2119 vss.n316 vss.n315 0.121289
R2120 vss.n316 vss.n298 0.121289
R2121 vss.n782 vss.n781 0.121289
R2122 vss.n781 vss.n780 0.121289
R2123 vss.n201 vss.n199 0.121289
R2124 vss.n287 vss.n199 0.121289
R2125 vss.n1478 vss.n56 0.121289
R2126 vss.n1473 vss.n56 0.121289
R2127 vss.n1473 vss.n1472 0.121289
R2128 vss.n1480 vss.n1479 0.121289
R2129 vss.n55 vss.n54 0.121289
R2130 vss.n54 vss.n10 0.121289
R2131 vss.n49 vss.n10 0.121289
R2132 vss.n49 vss.n48 0.121289
R2133 vss.n48 vss.n12 0.121289
R2134 vss.n43 vss.n12 0.121289
R2135 vss.n43 vss.n42 0.121289
R2136 vss.n42 vss.n41 0.121289
R2137 vss.n41 vss.n14 0.121289
R2138 vss.n35 vss.n14 0.121289
R2139 vss.n35 vss.n34 0.121289
R2140 vss.n34 vss.n33 0.121289
R2141 vss.n33 vss.n16 0.121289
R2142 vss.n27 vss.n16 0.121289
R2143 vss.n27 vss.n26 0.121289
R2144 vss.n26 vss.n25 0.121289
R2145 vss.n25 vss.n18 0.121289
R2146 vss.n19 vss.n18 0.121289
R2147 vss.n19 vss.n2 0.121289
R2148 vss.n177 vss.n160 0.121289
R2149 vss.n178 vss.n177 0.121289
R2150 vss.n153 vss.n90 0.121289
R2151 vss.n159 vss.n153 0.121289
R2152 vss.n370 vss.n366 0.121289
R2153 vss.n366 vss.n365 0.121289
R2154 vss.n765 vss.n299 0.121289
R2155 vss.n765 vss.n764 0.121289
R2156 vss.n415 vss.n403 0.121289
R2157 vss.n744 vss.n398 0.121289
R2158 vss.n416 vss.n398 0.121289
R2159 vss.n733 vss.n418 0.121289
R2160 vss.n733 vss.n732 0.121289
R2161 vss.n731 vss.n419 0.121289
R2162 vss.n751 vss.n390 0.121289
R2163 vss.n746 vss.n390 0.121289
R2164 vss.n280 vss.n182 0.121289
R2165 vss.n795 vss.n182 0.121289
R2166 vss.n1376 vss.n1375 0.121289
R2167 vss.n1375 vss.n1363 0.121289
R2168 vss.n1364 vss.n1363 0.121289
R2169 vss.n1377 vss.n1362 0.121289
R2170 vss.n1361 vss.n818 0.121289
R2171 vss.n1356 vss.n818 0.121289
R2172 vss.n1356 vss.n1355 0.121289
R2173 vss.n1355 vss.n1354 0.121289
R2174 vss.n1354 vss.n820 0.121289
R2175 vss.n1348 vss.n820 0.121289
R2176 vss.n1348 vss.n1347 0.121289
R2177 vss.n1347 vss.n1346 0.121289
R2178 vss.n1346 vss.n822 0.121289
R2179 vss.n1340 vss.n822 0.121289
R2180 vss.n1340 vss.n1339 0.121289
R2181 vss.n1339 vss.n1338 0.121289
R2182 vss.n1338 vss.n824 0.121289
R2183 vss.n1332 vss.n824 0.121289
R2184 vss.n1332 vss.n1331 0.121289
R2185 vss.n1331 vss.n1330 0.121289
R2186 vss.n1330 vss.n826 0.121289
R2187 vss.n1324 vss.n826 0.121289
R2188 vss.n1324 vss.n1323 0.121289
R2189 vss.n1304 vss.n1302 0.121289
R2190 vss.n1302 vss.n1299 0.121289
R2191 vss.n1299 vss.n1298 0.121289
R2192 vss.n1298 vss.n1295 0.121289
R2193 vss.n1295 vss.n1294 0.121289
R2194 vss.n1294 vss.n1291 0.121289
R2195 vss.n1291 vss.n1290 0.121289
R2196 vss.n1290 vss.n1287 0.121289
R2197 vss.n1287 vss.n830 0.121289
R2198 vss.n1318 vss.n830 0.121289
R2199 vss.n1306 vss.n1305 0.121289
R2200 vss.n1286 vss.n1285 0.121289
R2201 vss.n1285 vss.n861 0.121289
R2202 vss.n1280 vss.n861 0.121289
R2203 vss.n1059 vss.n949 0.121289
R2204 vss.n1059 vss.n1058 0.121289
R2205 vss.n986 vss.n977 0.121289
R2206 vss.n981 vss.n977 0.121289
R2207 vss.n1003 vss.n987 0.121289
R2208 vss.n1003 vss.n1002 0.121289
R2209 vss.n994 vss.n993 0.121289
R2210 vss.n994 vss.n989 0.121289
R2211 vss.n1000 vss.n989 0.121289
R2212 vss.n1441 vss.n1440 0.120962
R2213 vss.n1415 vss.n121 0.119721
R2214 vss.n1415 vss.n1414 0.119721
R2215 vss.n235 vss.n234 0.119721
R2216 vss.n245 vss.n235 0.119721
R2217 vss.n1245 vss.n864 0.119721
R2218 vss.n1277 vss.n864 0.119721
R2219 vss.n1185 vss.n1184 0.116268
R2220 vss.n624 vss.n623 0.106112
R2221 vss.n992 vss.n991 0.104479
R2222 vss.n171 vss.n170 0.100283
R2223 vss.n687 vss.n686 0.0994399
R2224 vss.n1194 vss.n1187 0.0942344
R2225 vss.n1319 vss.n1318 0.0928684
R2226 vss.n772 vss.n771 0.0923
R2227 vss.n1485 vss.n1484 0.0867105
R2228 vss.n609 vss.n608 0.084579
R2229 vss.n1472 vss.n1471 0.0839545
R2230 vss.n1367 vss.n1364 0.0839545
R2231 vss.n1280 vss.n1279 0.0839545
R2232 vss.n1322 vss.n1321 0.0828116
R2233 vss.n648 vss.n647 0.0824838
R2234 vss.n706 vss.n705 0.0824838
R2235 vss.n707 vss.n706 0.0824838
R2236 vss.n798 vss.n180 0.0817389
R2237 vss.n798 vss.n797 0.0817389
R2238 vss.n327 vss.n185 0.0817389
R2239 vss.n328 vss.n327 0.0817389
R2240 vss.n329 vss.n328 0.0817389
R2241 vss.n379 vss.n324 0.0817389
R2242 vss.n380 vss.n379 0.0817389
R2243 vss.n381 vss.n380 0.0817389
R2244 vss.n762 vss.n382 0.0817389
R2245 vss.n395 vss.n382 0.0817389
R2246 vss.n397 vss.n395 0.0817389
R2247 vss.n1196 vss.n1194 0.0814651
R2248 vss.n1184 vss.n1183 0.0807905
R2249 vss.n713 vss.n427 0.077759
R2250 vss.n966 vss.n962 0.076587
R2251 vss.n773 vss.n772 0.0739969
R2252 vss.n676 vss 0.0720663
R2253 vss.n815 vss.n813 0.0712322
R2254 vss.n632 vss.n631 0.0704647
R2255 vss.n754 vss.n753 0.0695
R2256 vss.n740 vss.n389 0.0685
R2257 vss.n740 vss.n739 0.0685
R2258 vss.n737 vss.n404 0.0685
R2259 vss.n726 vss.n404 0.0685
R2260 vss.n170 vss.n162 0.0664166
R2261 vss.n616 vss.n496 0.06425
R2262 vss.n611 vss.n496 0.06425
R2263 vss.n611 vss.n610 0.06425
R2264 vss.n583 vss.n506 0.06425
R2265 vss.n584 vss.n583 0.06425
R2266 vss.n587 vss.n584 0.06425
R2267 vss.n588 vss.n587 0.06425
R2268 vss.n591 vss.n588 0.06425
R2269 vss.n593 vss.n591 0.06425
R2270 vss.n771 vss.n300 0.0617
R2271 vss.n755 vss.n300 0.0617
R2272 vss.n755 vss.n754 0.0617
R2273 vss.n626 vss 0.0615976
R2274 vss.n609 vss.n506 0.059875
R2275 vss.n1413 vss.n122 0.0598265
R2276 vss.n244 vss.n243 0.0598265
R2277 vss.n1244 vss.n1243 0.0598265
R2278 vss.n1196 vss.n1195 0.0597258
R2279 vss.n1229 vss.n1222 0.0596781
R2280 vss.n1273 vss.n1272 0.0596781
R2281 vss.n113 vss.n107 0.0596781
R2282 vss.n224 vss.n82 0.0596781
R2283 vss.n1401 vss.n144 0.0572123
R2284 vss.n252 vss.n250 0.0572123
R2285 vss.n1057 vss.n1056 0.0542097
R2286 vss.n599 vss.n593 0.053625
R2287 vss.n1136 vss.n1110 0.0525435
R2288 vss.n1100 vss.n1074 0.0525435
R2289 vss.n564 vss.n563 0.0525312
R2290 vss.n354 vss.n288 0.0525312
R2291 vss.n920 vss.n919 0.0524302
R2292 vss vss.n961 0.0518423
R2293 vss.n752 vss.n751 0.0502368
R2294 vss.n1039 vss.n1026 0.0500277
R2295 vss.n1039 vss.n1038 0.0500277
R2296 vss.n622 vss.n491 0.0488158
R2297 vss.n1484 vss.n3 0.0488158
R2298 vss.n1008 vss.n1007 0.0487143
R2299 vss.n1195 vss.n1 0.0469516
R2300 vss.n1321 vss.n815 0.0466307
R2301 vss vss.n1186 0.0449398
R2302 vss.n706 vss.n434 0.0442727
R2303 vss.n692 vss.n444 0.0442727
R2304 vss.n1391 vss.n131 0.0428443
R2305 vss.n1222 vss.n872 0.0424178
R2306 vss.n1273 vss.n872 0.0424178
R2307 vss.n148 vss.n113 0.0424178
R2308 vss.n149 vss.n148 0.0424178
R2309 vss.n224 vss.n218 0.0424178
R2310 vss.n249 vss.n218 0.0424178
R2311 vss.n486 vss.n480 0.0422273
R2312 vss.n489 vss.n486 0.0422273
R2313 vss.n490 vss.n489 0.0422273
R2314 vss.n693 vss.n434 0.0422273
R2315 vss.n693 vss.n692 0.0422273
R2316 vss.n1470 vss.n1467 0.0422273
R2317 vss.n1460 vss.n1457 0.0422273
R2318 vss.n1457 vss.n1456 0.0422273
R2319 vss.n1453 vss.n1452 0.0422273
R2320 vss.n1368 vss.n100 0.0422273
R2321 vss.n1428 vss.n1427 0.0422273
R2322 vss.n1427 vss.n1426 0.0422273
R2323 vss.n1421 vss.n109 0.0422273
R2324 vss.n881 vss.n863 0.0422273
R2325 vss.n892 vss.n891 0.0422273
R2326 vss.n892 vss.n873 0.0422273
R2327 vss.n1271 vss.n874 0.0422273
R2328 vss.n1260 vss.n899 0.0422273
R2329 vss.n1255 vss.n899 0.0422273
R2330 vss.n1255 vss.n1254 0.0422273
R2331 vss.n1443 vss.n1442 0.0414091
R2332 vss.n1388 vss.n1387 0.0414091
R2333 vss.n677 vss.n676 0.0407439
R2334 vss.n1040 vss.n1039 0.0404194
R2335 vss.n1145 vss.n1110 0.040413
R2336 vss.n1163 vss.n1074 0.040413
R2337 vss.n556 vss.n555 0.0391719
R2338 vss.n363 vss.n361 0.0391719
R2339 vss vss.n920 0.0389394
R2340 vss.n555 vss.n554 0.0388607
R2341 vss.n1389 vss.n1388 0.0379754
R2342 vss.n626 vss.n625 0.0378171
R2343 vss.n625 vss.n455 0.0378171
R2344 vss.n665 vss.n664 0.0378171
R2345 vss.n666 vss.n665 0.0378171
R2346 vss.n667 vss.n666 0.0378171
R2347 vss.n678 vss.n677 0.0378171
R2348 vss.n649 vss.n648 0.037666
R2349 vss.n649 vss.n435 0.037666
R2350 vss.n705 vss.n435 0.037666
R2351 vss.n708 vss.n707 0.037666
R2352 vss.n708 vss.n425 0.037666
R2353 vss.n721 vss.n425 0.037666
R2354 vss.n1056 vss.n951 0.0375161
R2355 vss.n1051 vss.n951 0.0375161
R2356 vss.n1051 vss.n1050 0.0375161
R2357 vss.n1050 vss.n1048 0.0375161
R2358 vss.n1048 vss.n1044 0.0375161
R2359 vss.n1044 vss.n1043 0.0375161
R2360 vss.n1043 vss.n1040 0.0375161
R2361 vss.n609 vss.n507 0.0372105
R2362 vss.n1153 vss 0.0368913
R2363 vss.n1171 vss 0.0368913
R2364 vss.n563 vss.n520 0.0363594
R2365 vss.n531 vss.n520 0.0363594
R2366 vss.n532 vss.n531 0.0363594
R2367 vss.n536 vss.n532 0.0363594
R2368 vss.n538 vss.n536 0.0363594
R2369 vss.n557 vss.n538 0.0363594
R2370 vss.n557 vss.n556 0.0363594
R2371 vss.n354 vss.n353 0.0363594
R2372 vss.n353 vss.n352 0.0363594
R2373 vss.n352 vss.n349 0.0363594
R2374 vss.n349 vss.n345 0.0363594
R2375 vss.n345 vss.n338 0.0363594
R2376 vss.n360 vss.n338 0.0363594
R2377 vss.n361 vss.n360 0.0363594
R2378 vss.n1453 vss.n82 0.0360909
R2379 vss.n109 vss.n107 0.0360909
R2380 vss.n1272 vss.n1271 0.0360909
R2381 vss.n1406 vss.n131 0.0351154
R2382 vss.n269 vss.n268 0.0351154
R2383 vss.n1234 vss.n920 0.0351154
R2384 vss.n634 vss.n632 0.0344545
R2385 vss.n1146 vss.n1109 0.0337609
R2386 vss.n1164 vss.n1073 0.0337609
R2387 vss.n701 vss.n700 0.0329382
R2388 vss.n685 vss.n684 0.0329382
R2389 vss.n139 vss.n138 0.0325979
R2390 vss.n143 vss.n142 0.0325979
R2391 vss.n1402 vss.n143 0.0325979
R2392 vss.n1400 vss.n147 0.0325979
R2393 vss.n242 vss.n236 0.0325979
R2394 vss.n237 vss.n217 0.0325979
R2395 vss.n253 vss.n217 0.0325979
R2396 vss.n251 vss.n214 0.0325979
R2397 vss.n1242 vss.n910 0.0325979
R2398 vss.n1221 vss.n1218 0.0325979
R2399 vss.n1230 vss.n1221 0.0325979
R2400 vss.n1228 vss.n1225 0.0325979
R2401 vss.n475 vss.n463 0.0324091
R2402 vss.n641 vss.n640 0.0324091
R2403 vss.n635 vss.n476 0.0324091
R2404 vss.n169 vss.n167 0.0323462
R2405 vss.n654 vss.n460 0.0313481
R2406 vss.n659 vss.n655 0.0313481
R2407 vss.n658 vss.n657 0.0313481
R2408 vss.n701 vss.n443 0.0313481
R2409 vss.n555 vss 0.0298607
R2410 vss.n1467 vss.n1466 0.0291364
R2411 vss.n78 vss.n70 0.0291364
R2412 vss.n1461 vss.n81 0.0291364
R2413 vss.n1434 vss.n100 0.0291364
R2414 vss.n1433 vss.n101 0.0291364
R2415 vss.n106 vss.n103 0.0291364
R2416 vss.n881 vss.n877 0.0291364
R2417 vss.n886 vss.n885 0.0291364
R2418 vss.n890 vss.n876 0.0291364
R2419 vss vss.n1487 0.029
R2420 vss.n714 vss.n713 0.0286928
R2421 vss.n673 vss.n427 0.0281506
R2422 vss.n1252 vss.n1251 0.0271119
R2423 vss.n1442 vss.n1441 0.0269232
R2424 vss.n647 vss.n646 0.0267348
R2425 vss.n1252 vss.n855 0.0266818
R2426 vss.n270 vss.n206 0.0259844
R2427 vss.n753 vss.n752 0.0258333
R2428 vss.n1452 vss.n83 0.0254545
R2429 vss.n1449 vss.n1448 0.0254545
R2430 vss.n1446 vss.n84 0.0254545
R2431 vss.n1421 vss.n1420 0.0254545
R2432 vss.n810 vss.n111 0.0254545
R2433 vss.n811 vss.n807 0.0254545
R2434 vss.n897 vss.n874 0.0254545
R2435 vss.n1266 vss.n1265 0.0254545
R2436 vss.n1261 vss.n898 0.0254545
R2437 vss.n1194 vss.n1193 0.0253684
R2438 vss.n431 vss.n430 0.025235
R2439 vss.n597 vss.n595 0.0251316
R2440 vss.n372 vss.n371 0.0250455
R2441 vss.n1401 vss.n1400 0.0247308
R2442 vss.n252 vss.n251 0.0247308
R2443 vss.n1229 vss.n1228 0.0247308
R2444 vss.n685 vss.n444 0.0246696
R2445 vss.n595 vss.n491 0.0241842
R2446 vss.n1109 vss.n1103 0.023587
R2447 vss.n1073 vss.n1067 0.023587
R2448 vss.n632 vss.n482 0.0233975
R2449 vss.n147 vss.n145 0.0228427
R2450 vss.n1409 vss.n130 0.0228427
R2451 vss.n1408 vss.n1407 0.0228427
R2452 vss.n214 vss.n212 0.0228427
R2453 vss.n262 vss.n261 0.0228427
R2454 vss.n263 vss.n207 0.0228427
R2455 vss.n1225 vss.n1223 0.0228427
R2456 vss.n1237 vss.n918 0.0228427
R2457 vss.n1236 vss.n1235 0.0228427
R2458 vss.n580 vss.n579 0.0223361
R2459 vss.n668 vss.n667 0.0217195
R2460 vss.n1441 vss.n89 0.0212692
R2461 vss.n1001 vss.n988 0.0209545
R2462 vss.n1024 vss.n961 0.0206745
R2463 vss.n1319 vss.n828 0.0206316
R2464 vss.n713 vss.n712 0.0205353
R2465 vss.n455 vss.n453 0.0202561
R2466 vss vss.n624 0.0198902
R2467 vss.n1026 vss.n1025 0.0193501
R2468 vss.n1038 vss.n1027 0.0193501
R2469 vss.n1030 vss.n1027 0.0193501
R2470 vss.n1250 vss.n902 0.0193501
R2471 vss.n1251 vss.n1250 0.0193501
R2472 vss.n664 vss.n453 0.018061
R2473 vss.n683 vss.n428 0.0179912
R2474 vss vss.n541 0.0177623
R2475 vss.n632 vss.n480 0.0176818
R2476 vss.n624 vss.n490 0.0176818
R2477 vss.n1152 vss.n1103 0.0173261
R2478 vss.n1170 vss.n1067 0.0173261
R2479 vss.n1449 vss.n83 0.0172727
R2480 vss.n1448 vss.n1446 0.0172727
R2481 vss.n1443 vss.n84 0.0172727
R2482 vss.n1420 vss.n111 0.0172727
R2483 vss.n811 vss.n810 0.0172727
R2484 vss.n1387 vss.n807 0.0172727
R2485 vss.n1266 vss.n897 0.0172727
R2486 vss.n1265 vss.n898 0.0172727
R2487 vss.n1261 vss.n1260 0.0172727
R2488 vss.n1001 vss.n1000 0.0171646
R2489 vss.n678 vss.n668 0.0165976
R2490 vss.n1025 vss.n1024 0.0164061
R2491 vss vss.n1152 0.0161522
R2492 vss vss.n1170 0.0161522
R2493 vss.n1254 vss.n1252 0.0160455
R2494 vss.n1017 vss.n967 0.0155852
R2495 vss.n1016 vss.n968 0.0155852
R2496 vss.n1011 vss.n963 0.0155852
R2497 vss.n542 vss.n540 0.0155492
R2498 vss.n553 vss.n540 0.0155492
R2499 vss.n578 vss.n513 0.0155492
R2500 vss.n579 vss.n578 0.0155492
R2501 vss.n1390 vss.n1389 0.0155492
R2502 vss.n684 vss.n683 0.015447
R2503 vss.n712 vss.n428 0.015447
R2504 vss.n1030 vss 0.0150996
R2505 vss.n229 vss.n88 0.0141811
R2506 vss.n229 vss.n206 0.0141811
R2507 vss.n277 vss.n205 0.0141811
R2508 vss.n362 vss.n190 0.0141811
R2509 vss.n775 vss.n774 0.0141811
R2510 vss vss.n277 0.0140469
R2511 vss.n541 vss.n131 0.0139262
R2512 vss.n279 vss.n189 0.0139128
R2513 vss.n1466 vss.n70 0.0135909
R2514 vss.n81 vss.n78 0.0135909
R2515 vss.n1461 vss.n1460 0.0135909
R2516 vss.n1434 vss.n1433 0.0135909
R2517 vss.n103 vss.n101 0.0135909
R2518 vss.n1428 vss.n106 0.0135909
R2519 vss.n885 vss.n877 0.0135909
R2520 vss.n886 vss.n876 0.0135909
R2521 vss.n891 vss.n890 0.0135909
R2522 vss.n270 vss.n269 0.0135104
R2523 vss.n1007 vss.n1006 0.0134262
R2524 vss.n647 vss.n463 0.0123636
R2525 vss.n363 vss.n362 0.0121692
R2526 vss.n542 vss 0.0121557
R2527 vss.n926 vss.n1 0.0116429
R2528 vss.n789 vss.n189 0.0116326
R2529 vss.n788 vss.n190 0.0116326
R2530 vss.n988 vss.n967 0.0114943
R2531 vss.n1017 vss.n1016 0.0114943
R2532 vss.n1011 vss.n968 0.0114943
R2533 vss vss.n513 0.0112705
R2534 vss.n599 vss.n598 0.011125
R2535 vss.n278 vss 0.0110961
R2536 vss.n335 vss.n194 0.0110961
R2537 vss.n334 vss.n333 0.0110961
R2538 vss.n775 vss.n297 0.0110961
R2539 vss.n220 vss.n215 0.0108879
R2540 vss.n371 vss.n194 0.0104255
R2541 vss.n641 vss.n475 0.0103182
R2542 vss.n640 vss.n476 0.0103182
R2543 vss.n635 vss.n634 0.0103182
R2544 vss.n145 vss.n130 0.0102552
R2545 vss.n1409 vss.n1408 0.0102552
R2546 vss.n1407 vss.n1406 0.0102552
R2547 vss.n261 vss.n212 0.0102552
R2548 vss.n263 vss.n262 0.0102552
R2549 vss.n268 vss.n207 0.0102552
R2550 vss.n1223 vss.n918 0.0102552
R2551 vss.n1237 vss.n1236 0.0102552
R2552 vss.n1235 vss.n1234 0.0102552
R2553 vss.n1442 vss.n87 0.0101572
R2554 vss.n1009 vss.n1008 0.0101429
R2555 vss.n700 vss.n444 0.00876855
R2556 vss vss.n1390 0.00861475
R2557 vss.n1402 vss.n1401 0.00836713
R2558 vss.n253 vss.n252 0.00836713
R2559 vss.n1230 vss.n1229 0.00836713
R2560 vss.n1441 vss.n88 0.00814531
R2561 vss.n138 vss.n122 0.00805245
R2562 vss.n243 vss.n242 0.00805245
R2563 vss.n1243 vss.n1242 0.00805245
R2564 vss.n161 vss.n160 0.00760526
R2565 vss.n1388 vss.n806 0.00758197
R2566 vss.n1366 vss.n121 0.00751299
R2567 vss.n234 vss.n69 0.00751299
R2568 vss.n1278 vss.n1277 0.00751299
R2569 vss.n1391 vss 0.00743443
R2570 vss.n142 vss.n139 0.00742308
R2571 vss.n237 vss.n236 0.00742308
R2572 vss.n1218 vss.n910 0.00742308
R2573 vss.n1146 vss.n1145 0.00715217
R2574 vss.n1164 vss.n1163 0.00715217
R2575 vss.n1456 vss.n82 0.00663636
R2576 vss.n1426 vss.n107 0.00663636
R2577 vss.n1272 vss.n873 0.00663636
R2578 vss.n600 vss.n599 0.00610656
R2579 vss.n185 vss.n181 0.00607522
R2580 vss.n168 vss.n87 0.00559687
R2581 vss.n600 vss.n580 0.00551639
R2582 vss.n610 vss.n609 0.004875
R2583 vss.n813 vss.n806 0.00404098
R2584 vss.n335 vss.n334 0.00358495
R2585 vss.n333 vss.n297 0.00358495
R2586 vss.n623 vss.n622 0.00334211
R2587 vss.n789 vss.n788 0.00304844
R2588 vss.n149 vss.n144 0.00296575
R2589 vss.n250 vss.n249 0.00296575
R2590 vss.n1471 vss.n1470 0.00295455
R2591 vss.n1368 vss.n1367 0.00295455
R2592 vss.n1279 vss.n863 0.00295455
R2593 vss.n372 vss.n363 0.00251192
R2594 vss.n554 vss.n553 0.00227049
R2595 vss.n631 vss.n460 0.00209011
R2596 vss.n655 vss.n654 0.00209011
R2597 vss.n659 vss.n658 0.00209011
R2598 vss.n657 vss.n443 0.00209011
R2599 vss.n1007 vss 0.00194966
R2600 vss.n919 vss.n902 0.00160883
R2601 vss vss.n673 0.00131325
R2602 vss.n269 vss.n205 0.00117064
R2603 vss.n279 vss.n278 0.000768256
R2604 vss.n774 vss.n773 0.000634128
R2605 vdd.t53 vdd.t21 933.037
R2606 vdd.t21 vdd.t23 834.822
R2607 vdd.t62 vdd.t64 715.827
R2608 vdd.t45 vdd.t65 594.059
R2609 vdd.n30 vdd.t38 501.8
R2610 vdd.n108 vdd.t39 501.8
R2611 vdd.t39 vdd 489.991
R2612 vdd.n33 vdd.t38 489.502
R2613 vdd.n31 vdd.t62 489.219
R2614 vdd.n38 vdd.t60 489.219
R2615 vdd.n68 vdd.t16 476.993
R2616 vdd.t64 vdd.n30 476.62
R2617 vdd.t65 vdd.n108 476.62
R2618 vdd.t60 vdd.n37 336.332
R2619 vdd.n62 vdd.n58 330.935
R2620 vdd.t18 vdd.n63 311.151
R2621 vdd.t16 vdd.t0 306.656
R2622 vdd.n50 vdd.n47 277.878
R2623 vdd.n44 vdd.t56 266.188
R2624 vdd.n110 vdd.n109 256.137
R2625 vdd.n35 vdd.t32 250.899
R2626 vdd.n41 vdd.t32 244.75
R2627 vdd.n52 vdd.t25 238.31
R2628 vdd.n55 vdd.t66 238.31
R2629 vdd.t28 vdd.n56 238.31
R2630 vdd.n67 vdd.t49 238.31
R2631 vdd.t58 vdd.n45 215.827
R2632 vdd.t33 vdd.t58 215.827
R2633 vdd.t30 vdd.t41 201.44
R2634 vdd.t25 vdd.n51 197.843
R2635 vdd.t47 vdd.t2 191.548
R2636 vdd.n46 vdd.t26 178.958
R2637 vdd.n57 vdd.t55 178.059
R2638 vdd.t43 vdd.n50 160.072
R2639 vdd.n51 vdd.t34 160.072
R2640 vdd.t40 vdd.t33 142.087
R2641 vdd.t20 vdd.t36 131.296
R2642 vdd.t68 vdd.t18 126.799
R2643 vdd.n66 vdd.n64 126.799
R2644 vdd.t49 vdd.n66 124.102
R2645 vdd.n109 vdd.t45 117.007
R2646 vdd.n64 vdd.t68 111.511
R2647 vdd.n37 vdd.t20 107.014
R2648 vdd.t36 vdd.n35 107.014
R2649 vdd.t41 vdd.t28 102.519
R2650 vdd.n56 vdd.n55 90.8278
R2651 vdd.t34 vdd.t43 78.2379
R2652 vdd.t0 vdd.n67 69.2451
R2653 vdd.n12 vdd.n11 62.0058
R2654 vdd.n151 vdd.n150 62.0058
R2655 vdd.n99 vdd.n98 62.0058
R2656 vdd.n109 vdd.t53 60.2684
R2657 vdd.n58 vdd.n57 60.2523
R2658 vdd.t26 vdd.t40 59.353
R2659 vdd.n3 vdd.n2 54.711
R2660 vdd.n140 vdd.n139 54.711
R2661 vdd.n130 vdd.n93 54.711
R2662 vdd.n114 vdd.n106 54.5452
R2663 vdd.n115 vdd.n114 54.5452
R2664 vdd.t55 vdd.t30 53.9573
R2665 vdd.n47 vdd.n46 53.0581
R2666 vdd.n116 vdd.n115 48.3037
R2667 vdd.t2 vdd.n62 46.7631
R2668 vdd.n63 vdd.t47 46.7631
R2669 vdd.n7 vdd.n6 44.4321
R2670 vdd.n21 vdd.n7 44.4321
R2671 vdd.n144 vdd.n143 44.4321
R2672 vdd.n160 vdd.n144 44.4321
R2673 vdd.n128 vdd.n94 44.4321
R2674 vdd.n129 vdd.n128 44.4321
R2675 vdd.n14 vdd.n13 44.1177
R2676 vdd.n153 vdd.n152 44.1177
R2677 vdd.n122 vdd.n121 41.0086
R2678 vdd.n14 vdd.n5 31.6537
R2679 vdd.n153 vdd.n142 31.6537
R2680 vdd.n123 vdd.n122 31.6537
R2681 vdd.n13 vdd.n12 29.9841
R2682 vdd.n152 vdd.n151 29.9841
R2683 vdd.n120 vdd.n98 29.9841
R2684 vdd.n6 vdd.n2 29.5043
R2685 vdd.n143 vdd.n139 29.5043
R2686 vdd.n130 vdd.n129 29.5043
R2687 vdd.n106 vdd.n97 28.5602
R2688 vdd.n166 vdd.t8 26.892
R2689 vdd.n146 vdd.t6 24.3938
R2690 vdd.n23 vdd.n22 23.3768
R2691 vdd.n162 vdd.n161 23.3768
R2692 vdd.n96 vdd.n92 23.3768
R2693 vdd.n45 vdd.n44 22.4825
R2694 vdd.n34 vdd.n33 20.4586
R2695 vdd.n89 vdd.n41 20.2319
R2696 vdd.n11 vdd.n3 19.8952
R2697 vdd.n150 vdd.n140 19.8952
R2698 vdd.n99 vdd.n93 19.8952
R2699 vdd vdd.n146 19.301
R2700 vdd.n170 vdd.n169 19.1102
R2701 vdd.n89 vdd 18.6524
R2702 vdd.n29 vdd.n28 18.5371
R2703 vdd.n167 vdd.n166 18.4336
R2704 vdd.n28 vdd.n27 18.3436
R2705 vdd.n169 vdd.n168 18.3436
R2706 vdd.n135 vdd.n134 18.3436
R2707 vdd.n136 vdd.n135 18.3166
R2708 vdd.n27 vdd.t13 13.1071
R2709 vdd.n168 vdd.t11 13.1071
R2710 vdd.n146 vdd.t7 13.1071
R2711 vdd.n134 vdd.t15 13.1071
R2712 vdd.n32 vdd.n30 12.8823
R2713 vdd.n108 vdd.n107 12.8823
R2714 vdd.n69 vdd.n67 12.8823
R2715 vdd.n72 vdd.n64 12.8823
R2716 vdd.n76 vdd.n58 12.8823
R2717 vdd.n85 vdd.n46 12.8823
R2718 vdd.n77 vdd.n57 12.8823
R2719 vdd.n84 vdd.n47 12.8823
R2720 vdd vdd.n52 12.8823
R2721 vdd.n40 vdd.n35 12.8823
R2722 vdd.n45 vdd.n43 12.6005
R2723 vdd.n51 vdd.n49 12.6005
R2724 vdd.n55 vdd.n53 12.6005
R2725 vdd.n63 vdd.n60 12.6005
R2726 vdd.n66 vdd.n65 12.6005
R2727 vdd.n44 vdd.n42 12.6005
R2728 vdd.n50 vdd.n48 12.6005
R2729 vdd.n56 vdd.n54 12.6005
R2730 vdd.n62 vdd.n59 12.6005
R2731 vdd.n37 vdd.n36 12.6005
R2732 vdd.n166 vdd.t9 10.8823
R2733 vdd.n22 vdd.n4 10.8334
R2734 vdd.n161 vdd.n141 10.8334
R2735 vdd.n100 vdd.n96 10.8334
R2736 vdd.n10 vdd.n4 9.75782
R2737 vdd.n24 vdd.n23 9.75782
R2738 vdd.n149 vdd.n141 9.75782
R2739 vdd.n163 vdd.n162 9.75782
R2740 vdd.n131 vdd.n92 9.75782
R2741 vdd.n101 vdd.n100 9.75782
R2742 vdd vdd.t50 9.21665
R2743 vdd.n16 vdd.t5 8.94208
R2744 vdd.n17 vdd.t4 8.94208
R2745 vdd.n155 vdd.t52 8.94208
R2746 vdd.n156 vdd.t51 8.94208
R2747 vdd.n105 vdd.t22 8.94208
R2748 vdd.n126 vdd.t24 8.94208
R2749 vdd.n68 vdd.t17 8.42234
R2750 vdd.n70 vdd.t1 8.42234
R2751 vdd.n78 vdd.t31 8.42234
R2752 vdd.n79 vdd.t42 8.42234
R2753 vdd.n86 vdd.t27 8.42234
R2754 vdd.n31 vdd.t63 8.31339
R2755 vdd.n110 vdd.t46 8.31339
R2756 vdd.n59 vdd.t48 8.31339
R2757 vdd.n54 vdd.t29 8.31339
R2758 vdd.n48 vdd.t35 8.31339
R2759 vdd.n42 vdd.t59 8.31339
R2760 vdd.n36 vdd.t37 8.31339
R2761 vdd.n38 vdd.t61 8.31339
R2762 vdd.n65 vdd.t69 8.30475
R2763 vdd.n60 vdd.t3 8.30475
R2764 vdd.n53 vdd.t67 8.30475
R2765 vdd.n49 vdd.t44 8.30475
R2766 vdd.n43 vdd.t57 8.30475
R2767 vdd.n61 vdd.t19 8.1405
R2768 vdd.n23 vdd.n3 6.79787
R2769 vdd.n162 vdd.n140 6.79787
R2770 vdd.n93 vdd.n92 6.79787
R2771 vdd.n116 vdd.n97 4.97256
R2772 vdd.n22 vdd.n21 3.64787
R2773 vdd.n161 vdd.n160 3.64787
R2774 vdd.n96 vdd.n94 3.64787
R2775 vdd.n118 vdd.t54 3.52948
R2776 vdd.n121 vdd.n120 3.23339
R2777 vdd.n11 vdd.n4 3.1505
R2778 vdd.n150 vdd.n141 3.1505
R2779 vdd.n100 vdd.n99 3.1505
R2780 vdd.n27 vdd.t12 2.24244
R2781 vdd.n168 vdd.t10 2.24244
R2782 vdd.n134 vdd.t14 2.24244
R2783 vdd.n13 vdd.n8 2.1005
R2784 vdd.n21 vdd.n20 2.1005
R2785 vdd.n20 vdd.n5 2.1005
R2786 vdd.n6 vdd.n0 2.1005
R2787 vdd.n152 vdd.n145 2.1005
R2788 vdd.n160 vdd.n159 2.1005
R2789 vdd.n159 vdd.n142 2.1005
R2790 vdd.n143 vdd.n137 2.1005
R2791 vdd.n120 vdd.n119 2.1005
R2792 vdd.n129 vdd.n90 2.1005
R2793 vdd.n124 vdd.n123 2.1005
R2794 vdd.n124 vdd.n94 2.1005
R2795 vdd.t66 vdd.n52 1.79906
R2796 vdd.n22 vdd.n5 1.69074
R2797 vdd.n161 vdd.n142 1.69074
R2798 vdd.n123 vdd.n96 1.69074
R2799 vdd.n15 vdd.n14 1.5755
R2800 vdd.n18 vdd.n7 1.5755
R2801 vdd.n25 vdd.n24 1.5755
R2802 vdd.n10 vdd.n9 1.5755
R2803 vdd.n154 vdd.n153 1.5755
R2804 vdd.n157 vdd.n144 1.5755
R2805 vdd.n149 vdd.n148 1.5755
R2806 vdd.n164 vdd.n163 1.5755
R2807 vdd.n111 vdd.n106 1.5755
R2808 vdd.n115 vdd.n104 1.5755
R2809 vdd.n128 vdd.n127 1.5755
R2810 vdd.n122 vdd.n95 1.5755
R2811 vdd.n132 vdd.n131 1.5755
R2812 vdd.n102 vdd.n101 1.5755
R2813 vdd.n12 vdd.n10 1.46026
R2814 vdd.n24 vdd.n2 1.46026
R2815 vdd.n151 vdd.n149 1.46026
R2816 vdd.n163 vdd.n139 1.46026
R2817 vdd.n131 vdd.n130 1.46026
R2818 vdd.n101 vdd.n98 1.46026
R2819 vdd.n32 vdd.n31 1.30857
R2820 vdd.n136 vdd.n89 1.286
R2821 vdd.n117 vdd.n116 1.05197
R2822 vdd.n114 vdd.n113 1.0505
R2823 vdd.n34 vdd.n29 0.922
R2824 vdd.n113 vdd.n104 0.779711
R2825 vdd.n112 vdd.n107 0.643822
R2826 vdd.n118 vdd.n104 0.622211
R2827 vdd.n15 vdd.n8 0.607567
R2828 vdd.n154 vdd.n145 0.607567
R2829 vdd.n39 vdd.n38 0.567196
R2830 vdd.n147 vdd 0.566593
R2831 vdd.n170 vdd.n136 0.5505
R2832 vdd.n121 vdd.n97 0.538578
R2833 vdd.n113 vdd.n112 0.512741
R2834 vdd.n28 vdd 0.498918
R2835 vdd.n135 vdd 0.498918
R2836 vdd.n33 vdd 0.491
R2837 vdd.n17 vdd.n0 0.48464
R2838 vdd.n156 vdd.n137 0.48464
R2839 vdd.n126 vdd.n90 0.48226
R2840 vdd vdd.n170 0.422
R2841 vdd.n61 vdd 0.395064
R2842 vdd.n9 vdd.n8 0.392291
R2843 vdd.n112 vdd.n110 0.309149
R2844 vdd vdd.n34 0.307
R2845 vdd.n26 vdd.n0 0.285895
R2846 vdd.n147 vdd.n145 0.285895
R2847 vdd.n165 vdd.n137 0.285895
R2848 vdd.n133 vdd.n90 0.285895
R2849 vdd.n19 vdd.n18 0.27928
R2850 vdd.n158 vdd.n157 0.27928
R2851 vdd.n127 vdd.n125 0.275922
R2852 vdd.n125 vdd.n95 0.275922
R2853 vdd.n87 vdd 0.263188
R2854 vdd.n73 vdd.n61 0.26172
R2855 vdd.n75 vdd.n59 0.261195
R2856 vdd.n80 vdd.n54 0.261195
R2857 vdd.n83 vdd.n48 0.261195
R2858 vdd.n88 vdd.n42 0.261195
R2859 vdd.n39 vdd.n36 0.261195
R2860 vdd.n169 vdd 0.247811
R2861 vdd.n41 vdd 0.24575
R2862 vdd.n71 vdd.n65 0.234974
R2863 vdd.n74 vdd.n60 0.234974
R2864 vdd.n81 vdd.n53 0.234974
R2865 vdd.n82 vdd.n49 0.234974
R2866 vdd.n87 vdd.n43 0.234974
R2867 vdd.n40 vdd.n39 0.218188
R2868 vdd.n71 vdd.n70 0.2075
R2869 vdd.n76 vdd.n75 0.205813
R2870 vdd.n84 vdd.n83 0.172625
R2871 vdd.n117 vdd.n105 0.165429
R2872 vdd.n19 vdd.n16 0.156354
R2873 vdd.n158 vdd.n155 0.156354
R2874 vdd vdd.n82 0.150688
R2875 vdd vdd.n81 0.150688
R2876 vdd vdd.n74 0.150688
R2877 vdd.n73 vdd 0.147312
R2878 vdd.n103 vdd.n102 0.138889
R2879 vdd vdd.n79 0.137188
R2880 vdd.n25 vdd.n1 0.136775
R2881 vdd.n9 vdd.n1 0.136775
R2882 vdd.n102 vdd.n91 0.136775
R2883 vdd.n132 vdd.n91 0.136775
R2884 vdd vdd.n88 0.134938
R2885 vdd.n69 vdd 0.132125
R2886 vdd.n79 vdd 0.127063
R2887 vdd.n74 vdd.n73 0.1265
R2888 vdd.n16 vdd.n15 0.123427
R2889 vdd.n18 vdd.n17 0.123427
R2890 vdd.n155 vdd.n154 0.123427
R2891 vdd.n157 vdd.n156 0.123427
R2892 vdd vdd.n32 0.122
R2893 vdd vdd.n107 0.122
R2894 vdd.n127 vdd.n126 0.121946
R2895 vdd.n105 vdd.n95 0.121946
R2896 vdd.n111 vdd.n103 0.117332
R2897 vdd.n125 vdd.n124 0.107
R2898 vdd.n26 vdd.n25 0.106897
R2899 vdd.n133 vdd.n132 0.106897
R2900 vdd.n20 vdd.n19 0.106625
R2901 vdd.n159 vdd.n158 0.106625
R2902 vdd vdd.n26 0.106221
R2903 vdd vdd.n133 0.106221
R2904 vdd.n164 vdd.n138 0.103436
R2905 vdd.n148 vdd.n138 0.103436
R2906 vdd vdd.n86 0.101187
R2907 vdd.n83 vdd 0.101187
R2908 vdd vdd.n78 0.101187
R2909 vdd vdd.n68 0.101187
R2910 vdd.n20 vdd.n1 0.090875
R2911 vdd.n159 vdd.n138 0.090875
R2912 vdd.n124 vdd.n91 0.090875
R2913 vdd.n29 vdd 0.0905
R2914 vdd.n78 vdd.n77 0.082625
R2915 vdd vdd.n167 0.0825588
R2916 vdd.n165 vdd.n164 0.080867
R2917 vdd.n148 vdd.n147 0.080867
R2918 vdd vdd.n165 0.0748848
R2919 vdd vdd.n72 0.071375
R2920 vdd.n72 vdd 0.06125
R2921 vdd vdd.n40 0.06125
R2922 vdd.n81 vdd.n80 0.055625
R2923 vdd.n119 vdd.n118 0.0534573
R2924 vdd.n86 vdd.n85 0.0494375
R2925 vdd.n119 vdd.n103 0.0460488
R2926 vdd.n77 vdd.n76 0.0381875
R2927 vdd.n85 vdd.n84 0.0336875
R2928 vdd.n75 vdd 0.0303125
R2929 vdd.n82 vdd 0.0280625
R2930 vdd.n70 vdd.n69 0.0201875
R2931 vdd vdd.n71 0.0190625
R2932 vdd.n88 vdd.n87 0.01625
R2933 vdd.n80 vdd 0.0156875
R2934 vdd.n112 vdd.n111 0.00329503
R2935 vdd.n167 vdd 0.00201261
R2936 vdd.n118 vdd.n117 0.00187113
R2937 v_rew v_rew.t3 37.2214
R2938 v_rew.n0 v_rew.t0 32.5076
R2939 v_rew.n1 v_rew.t2 28.3362
R2940 v_rew.n2 v_rew.t1 28.3362
R2941 v_rew.n2 v_rew.n1 11.0961
R2942 v_rew.n1 v_rew 5.4005
R2943 v_rew.n0 v_rew 4.71875
R2944 v_rew v_rew.n0 0.104711
R2945 v_rew v_rew.n2 0.102342
R2946 phi_fire.n0 phi_fire.t13 41.9396
R2947 phi_fire.n6 phi_fire.t5 41.9396
R2948 phi_fire.n3 phi_fire.t8 39.4319
R2949 phi_fire.n5 phi_fire.t15 37.4396
R2950 phi_fire.n9 phi_fire.t14 37.4396
R2951 phi_fire.n2 phi_fire.t9 34.4873
R2952 phi_fire.n11 phi_fire.t4 33.5205
R2953 phi_fire.n0 phi_fire.t16 32.5076
R2954 phi_fire.n4 phi_fire.t2 32.5076
R2955 phi_fire.n8 phi_fire.t12 32.5076
R2956 phi_fire.n6 phi_fire.t3 32.5076
R2957 phi_fire phi_fire.t7 28.457
R2958 phi_fire.n1 phi_fire.t6 28.3362
R2959 phi_fire.n3 phi_fire.t11 28.3362
R2960 phi_fire.n7 phi_fire.t10 28.3362
R2961 phi_fire.n14 phi_fire 12.9706
R2962 phi_fire.n10 phi_fire.n9 9.9725
R2963 phi_fire phi_fire.n13 9.2525
R2964 phi_fire phi_fire.t1 9.04888
R2965 phi_fire.n12 phi_fire.n11 9.0005
R2966 phi_fire.n14 phi_fire.t0 8.1405
R2967 phi_fire.n12 phi_fire.n5 6.15087
R2968 phi_fire.n10 phi_fire.n7 5.63162
R2969 phi_fire.n2 phi_fire.n1 4.94505
R2970 phi_fire.n5 phi_fire.n4 4.5005
R2971 phi_fire.n9 phi_fire.n8 4.5005
R2972 phi_fire.n13 phi_fire.n12 4.5005
R2973 phi_fire phi_fire.n14 0.332129
R2974 phi_fire.n13 phi_fire.n2 0.321125
R2975 phi_fire.n11 phi_fire.n10 0.255071
R2976 phi_fire phi_fire.n0 0.104711
R2977 phi_fire.n4 phi_fire 0.104711
R2978 phi_fire phi_fire.n6 0.104711
R2979 phi_fire.n1 phi_fire 0.102342
R2980 phi_fire phi_fire.n3 0.102342
R2981 phi_fire.n7 phi_fire 0.102342
R2982 phi_fire.n8 phi_fire 0.0857632
R2983 vmem vmem.t11 20.2482
R2984 vmem.n2 vmem.t4 16.4806
R2985 vmem.n2 vmem.n1 14.1316
R2986 vmem.n4 vmem.t3 13.1366
R2987 vmem.n7 vmem.n6 9.716
R2988 vmem.n5 vmem.n4 9.63725
R2989 vmem vmem.t5 9.17794
R2990 vmem vmem.t0 9.14522
R2991 vmem.n8 vmem.n7 9.0005
R2992 vmem.n0 vmem.t7 8.8205
R2993 vmem.n1 vmem.t9 8.8205
R2994 vmem vmem.t8 8.57004
R2995 vmem vmem.t10 8.53506
R2996 vmem.n8 vmem.t6 8.1405
R2997 vmem.n6 vmem.t1 8.1405
R2998 vmem.n3 vmem.n0 5.47925
R2999 vmem.n4 vmem.t2 4.99592
R3000 vmem vmem.n3 4.78962
R3001 vmem.n7 vmem.n5 2.507
R3002 vmem.n5 vmem 2.33487
R3003 vmem.n3 vmem.n2 0.818375
R3004 vmem vmem.n8 0.427318
R3005 vmem.n0 vmem 0.394944
R3006 vmem.n6 vmem 0.394591
R3007 vmem.n1 vmem 0.323598
R3008 vmem.n4 vmem 0.136625
R3009 vin.n0 vin.t4 59.6219
R3010 vin vin.t1 21.3485
R3011 vin.n3 vin.n2 18.652
R3012 vin.n1 vin.n0 18.5261
R3013 vin.n1 vin 12.01
R3014 vin.n3 vin.t2 8.8205
R3015 vin vin.t0 8.54078
R3016 vin vin.n3 0.38923
R3017 vin.n2 vin.t3 0.0455
R3018 vin.n2 vin.n1 0.0305
R3019 vin.n0 vin 0.003875
R3020 vout.n0 vout.t1 9.57203
R3021 vout vout.t2 9.21093
R3022 vout.n0 vout.t3 8.1405
R3023 vout.n2 vout.t0 8.1405
R3024 vout.n1 vout.n0 4.84475
R3025 vout.n2 vout.n1 4.5005
R3026 vout.n1 vout 0.856625
R3027 vout vout.n2 0.399071
C0 a_3544_2068# vspike 0.5989f
C1 v_rew phaseUpulse_0.phi_1 0.007f
C2 a_8075_6021# ota_1stage$2_0.vp 0.69632f
C3 a_2248_2068# vspike 0.59888f
C4 phaseUpulse_0.conmutator_0.out vspike 0.15135f
C5 a_2248_2068# a_3544_2068# 0.00376f
C6 v_rew phaseUpulse_0.vspike_down 0.00424f
C7 v_rew a_n872_2246# 0.79579f
C8 v_ref phaseUpulse_0.phi_2 0.02285f
C9 v_rew v_th 0.00409f
C10 phaseUpulse_0.phi_1 v_th 0.2582f
C11 a_n1388_602# phaseUpulse_0.monostable_0.not$1_3.in 0.00369f
C12 phaseUpulse_0.vspike_down a_n872_2246# 0
C13 phaseUpulse_0.monostable_0.not$1_1.in a_952_2068# 0.0012f
C14 phaseUpulse_0.monostable_0.nand$1_0.Z vspike 0.00176f
C15 a_n872_2246# v_th 0
C16 phaseUpulse_0.vspike_down v_th 0.40155f
C17 vdd phaseUpulse_0.phi_2 0.69232f
C18 phaseUpulse_0.vspike_down a_2328_3444# 0
C19 a_1251_5604# phaseUpulse_0.vspike_down 0.09495f
C20 a_1251_5604# v_th 0.00255f
C21 a_2328_3444# v_th 0.04862f
C22 v_rew phaseUpulse_0.vspike_up 0.35339f
C23 a_4045_6672# v_th 0
C24 a_8827_1078# phi_fire 0.94674f
C25 a_8811_n132# phi_fire 0.54852f
C26 vmem ota_1stage$2_0.vp 0.12636f
C27 a_6854_3116# vmem 0.03683f
C28 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_1 0.36261f
C29 phaseUpulse_0.vspike_up phaseUpulse_0.vspike_down 0.3677f
C30 phaseUpulse_0.vneg phaseUpulse_0.phi_1 0.33933f
C31 v_rew phaseUpulse_0.vneg 0.1251f
C32 phaseUpulse_0.vspike_up a_n872_2246# 0.08242f
C33 a_8827_1078# conmutator$1_2.out 0.75454f
C34 vout v_ref 0.1593f
C35 phaseUpulse_0.vspike_up v_th 0.03275f
C36 a_8811_n132# conmutator$1_2.out 0.0061f
C37 a_3790_3312# phi_fire 0.00627f
C38 a_6164_1900# vmem 0.1629f
C39 phaseUpulse_0.vspike_up a_1251_5604# 0.06422f
C40 phaseUpulse_0.vneg a_n872_2246# 0.02206f
C41 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.monostable_0.not$1_3.in 0.07366f
C42 phaseUpulse_0.monostable_0.not$1_0.in v_th 0.00666f
C43 phaseUpulse_0.vneg v_th 0.46093f
C44 phaseUpulse_0.monostable_0.nand$1_1.Z v_rew 0.02831f
C45 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.phi_1 0.00153f
C46 v_ref phi_fire 1.36814f
C47 a_8190_3623# vmem 1.01491f
C48 vout vdd 0.31925f
C49 conmutator$1_2.out v_ref 0.15117f
C50 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.phi_1 0
C51 a_9352_5200# vmem 0.50178f
C52 a_7562_3851# vmem 0.01101f
C53 phaseUpulse_0.monostable_0.nand$1_1.Z v_th 0.02529f
C54 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.vrefrac 0
C55 vdd phi_fire 3.89421f
C56 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.phi_2 0.04761f
C57 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vspike_down 0.07196f
C58 a_1078_602# phaseUpulse_0.monostable_0.nand$1_0.Z 0.04857f
C59 vmem vspike 0.09386f
C60 phaseUpulse_0.vspike_up phaseUpulse_0.vneg 0.04283f
C61 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_int 0
C62 conmutator$1_2.out vdd 0.4963f
C63 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn v_th 0.19924f
C64 v_ref phaseUpulse_0.phi_1 0.00326f
C65 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn a_2328_3444# 0.02667f
C66 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.vneg 0.004f
C67 a_3790_3312# v_th 0.00357f
C68 a_3544_1172# vdd 0.05888f
C69 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vspike_up 0.00609f
C70 v_rew ota_1stage$2_0.vout 0.07589f
C71 v_ref phaseUpulse_0.vspike_down 0
C72 a_3790_3312# a_2328_3444# 0.04633f
C73 vin phi_fire 0.28319f
C74 phaseUpulse_0.monostable_0.not$1_1.in vspike 0.00276f
C75 v_ref v_th 1.11094f
C76 vdd phaseUpulse_0.phi_1 1.6851f
C77 v_rew vdd 1.18265f
C78 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vspike_up 0
C79 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vneg 0.3112f
C80 phaseUpulse_0.vspike_down ota_1stage$2_0.vout 0.01354f
C81 a_n872_2246# ota_1stage$2_0.vout 0.00619f
C82 conmutator$1_2.out vin 0.79779f
C83 v_ref a_2328_3444# 0.01813f
C84 ota_1stage$2_0.vout v_th 0.02781f
C85 v_ref a_4045_6672# 0.00256f
C86 vdd phaseUpulse_0.vspike_down 0.1771f
C87 vdd a_n872_2246# 0.75706f
C88 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vneg 0.02731f
C89 a_1251_5604# ota_1stage$2_0.vout 0.01274f
C90 vdd v_th 1.00446f
C91 phaseUpulse_0.vrefrac phaseUpulse_0.phi_2 0.08553f
C92 a_2521_8244# v_th 0.00819f
C93 ota_1stage$2_0.vout a_4045_6672# 0
C94 vdd a_1251_5604# 0.00936f
C95 vdd a_2328_3444# 0.06355f
C96 a_8075_6021# vmem 0.08273f
C97 vdd a_4045_6672# 0.61031f
C98 phaseUpulse_0.phi_2 phaseUpulse_0.phi_int 0.25422f
C99 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.monostable_0.nand$1_0.Z 0.47226f
C100 a_2266_4884# phaseUpulse_0.phi_2 0
C101 a_2521_8244# a_4045_6672# 0.00553f
C102 phaseUpulse_0.vspike_up ota_1stage$2_0.vout 0.39904f
C103 vdd phaseUpulse_0.vspike_up 0.38521f
C104 a_8811_n132# a_8827_1078# 0
C105 vin v_th 0.04911f
C106 phaseUpulse_0.vneg ota_1stage$2_0.vout 0.20334f
C107 a_952_2068# phaseUpulse_0.phi_1 0.52142f
C108 v_rew a_952_2068# 0.00313f
C109 phaseUpulse_0.monostable_0.not$1_0.in vdd 0.60484f
C110 phaseUpulse_0.phi_2 vspike 0.27648f
C111 a_3790_3312# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0
C112 vdd phaseUpulse_0.vneg 0.80986f
C113 a_3544_2068# phaseUpulse_0.phi_2 0.0077f
C114 a_952_2068# a_n872_2246# 0.00376f
C115 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.phi_1 0.03454f
C116 a_952_2068# v_th 0.01009f
C117 phaseUpulse_0.monostable_0.nand$1_1.Z ota_1stage$2_0.vout 0.03281f
C118 a_8827_1078# v_ref 0.47663f
C119 a_1078_602# phaseUpulse_0.monostable_0.not$1_1.in 0.00369f
C120 a_2248_2068# phaseUpulse_0.phi_2 0.49862f
C121 ota_1stage$2_0.vp phi_fire 0.58514f
C122 a_6854_3116# phi_fire 0.02296f
C123 phaseUpulse_0.monostable_0.nand$1_1.Z vdd 0.41173f
C124 phaseUpulse_0.vspike_down phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0
C125 v_ref a_3790_3312# 0.26016f
C126 conmutator$1_2.out a_6854_3116# 0.00747f
C127 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp v_th 0.01894f
C128 vout a_8190_3623# 0.0164f
C129 a_6164_1900# phi_fire 0.06015f
C130 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn vdd 0.00279f
C131 a_1251_5604# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0
C132 a_8827_1078# vdd 0.28491f
C133 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp a_2328_3444# 0.09152f
C134 a_8811_n132# vdd 0.27677f
C135 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_2 0.00237f
C136 conmutator$1_2.out a_6164_1900# 0.03605f
C137 phaseUpulse_0.phi_int phi_fire 0.40552f
C138 v_rew phaseUpulse_0.monostable_0.not$1_3.in 0.0052f
C139 vout a_9352_5200# 0.69632f
C140 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.phi_1 0.00862f
C141 a_8190_3623# phi_fire 0.17771f
C142 a_3790_3312# vdd 0.58904f
C143 conmutator$1_2.out phaseUpulse_0.phi_int 0
C144 conmutator$1_2.out a_8190_3623# 0.00161f
C145 phaseUpulse_0.monostable_0.not$1_0.in a_952_2068# 0
C146 phaseUpulse_0.monostable_0.not$1_3.in a_n872_2246# 0
C147 a_9352_5200# phi_fire 0.86685f
C148 a_952_2068# phaseUpulse_0.vneg 0
C149 a_7562_3851# phi_fire 0.05873f
C150 v_ref vdd 0.88548f
C151 phaseUpulse_0.monostable_0.not$1_3.in v_th 0.07018f
C152 a_3544_1172# phaseUpulse_0.phi_int 0.04163f
C153 conmutator$1_2.out a_7562_3851# 0.00226f
C154 vspike phi_fire 0.11476f
C155 phaseUpulse_0.vrefrac phaseUpulse_0.phi_1 0.02211f
C156 a_8827_1078# vin 0.00869f
C157 a_8811_n132# vin 0.49018f
C158 a_3544_2068# phi_fire 0
C159 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.vneg 0.03166f
C160 vdd ota_1stage$2_0.vout 0.54064f
C161 v_th ota_1stage$2_0.vp 0.06191f
C162 conmutator$1_2.out vspike 0.06761f
C163 a_2521_8244# ota_1stage$2_0.vout 0.09327f
C164 phaseUpulse_0.phi_1 phaseUpulse_0.phi_int 0.05163f
C165 phaseUpulse_0.vrefrac phaseUpulse_0.vspike_down 0.00498f
C166 vdd a_2521_8244# 1.29114f
C167 v_th a_2583_6804# 0.04011f
C168 a_4045_6672# ota_1stage$2_0.vp 0.14528f
C169 phaseUpulse_0.vrefrac v_th 0.34655f
C170 a_3544_1172# vspike 0.00279f
C171 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.vspike_up 0
C172 a_3544_1172# a_3544_2068# 0
C173 a_2266_4884# phaseUpulse_0.vspike_down 0.01828f
C174 phaseUpulse_0.vrefrac a_2328_3444# 0.26447f
C175 vin v_ref 0.00374f
C176 a_4045_6672# a_2583_6804# 0.04633f
C177 a_2266_4884# v_th 0.2327f
C178 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.30977f
C179 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.vneg 0.42522f
C180 phaseUpulse_0.phi_1 vspike 0.48921f
C181 a_2328_3444# phaseUpulse_0.phi_int 0
C182 a_2266_4884# a_2328_3444# 0.39545f
C183 a_3544_2068# phaseUpulse_0.phi_1 0
C184 vin vdd 0.99519f
C185 a_3790_3312# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.01725f
C186 a_2248_2068# phaseUpulse_0.phi_1 0.00836f
C187 phaseUpulse_0.phi_1 phaseUpulse_0.conmutator_0.out 0.1136f
C188 v_rew phaseUpulse_0.conmutator_0.out 0.75989f
C189 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.monostable_0.not$1_3.in 0.47242f
C190 vspike v_th 0.00729f
C191 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.vrefrac 0
C192 a_8075_6021# phi_fire 0.87224f
C193 v_ref phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.01944f
C194 phaseUpulse_0.vrefrac phaseUpulse_0.vneg 0.00243f
C195 a_2328_3444# vspike 0
C196 vdd a_952_2068# 0.28111f
C197 a_n872_2246# phaseUpulse_0.conmutator_0.out 0.83515f
C198 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_int 0
C199 phaseUpulse_0.conmutator_0.out v_th 0.07567f
C200 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_1 0.2402f
C201 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_2 0.01642f
C202 vdd phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.01485f
C203 phaseUpulse_0.vrefrac phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0.30977f
C204 phaseUpulse_0.monostable_0.nand$1_0.Z v_th 0.17131f
C205 a_8827_1078# a_6164_1900# 0.00737f
C206 phaseUpulse_0.monostable_0.not$1_0.in vspike 0
C207 vout vmem 0.15077f
C208 phaseUpulse_0.vspike_up phaseUpulse_0.conmutator_0.out 0.09025f
C209 v_ref ota_1stage$2_0.vp 0.27429f
C210 phaseUpulse_0.monostable_0.not$1_3.in ota_1stage$2_0.vout 0.01206f
C211 phaseUpulse_0.vrefrac a_3790_3312# 0.01646f
C212 a_2266_4884# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0.00259f
C213 v_ref a_6854_3116# 0
C214 a_8827_1078# a_8190_3623# 0
C215 phaseUpulse_0.monostable_0.not$1_0.in a_2248_2068# 0
C216 a_1078_602# phaseUpulse_0.phi_1 0.00569f
C217 vdd phaseUpulse_0.monostable_0.not$1_3.in 0.2263f
C218 phaseUpulse_0.vneg phaseUpulse_0.conmutator_0.out 0.10052f
C219 vmem phi_fire 2.73321f
C220 a_3790_3312# phaseUpulse_0.phi_int 0.00115f
C221 a_2266_4884# a_3790_3312# 0.00553f
C222 v_ref phaseUpulse_0.vrefrac 0.00382f
C223 v_ref a_6164_1900# 0.00178f
C224 vdd ota_1stage$2_0.vp 0.49682f
C225 conmutator$1_2.out vmem 0.26299f
C226 a_n1388_602# v_rew 0
C227 vdd a_6854_3116# 0.06522f
C228 v_ref phaseUpulse_0.phi_int 0.23227f
C229 ota_1stage$2_0.vout a_2583_6804# 0.21159f
C230 a_2521_8244# ota_1stage$2_0.vp 0.03015f
C231 v_ref a_2266_4884# 0.03173f
C232 a_1078_602# v_th 0.00317f
C233 v_ref a_8190_3623# 0.24721f
C234 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.nand$1_0.Z 0.30883f
C235 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.conmutator_0.out 0
C236 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.vneg 0.00153f
C237 a_952_2068# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.00331f
C238 vdd a_2583_6804# 0.06682f
C239 phaseUpulse_0.vrefrac vdd 0.31314f
C240 vdd a_6164_1900# 0.53169f
C241 a_3790_3312# vspike 0.00965f
C242 a_2521_8244# a_2583_6804# 0.40678f
C243 v_ref a_9352_5200# 0.19585f
C244 a_3790_3312# a_3544_2068# 0.00141f
C245 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn a_2248_2068# 0
C246 v_ref a_7562_3851# 0
C247 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.conmutator_0.out 0.00674f
C248 vdd phaseUpulse_0.phi_int 0.70343f
C249 a_2266_4884# vdd 1.28499f
C250 vdd a_8190_3623# 1.10527f
C251 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.monostable_0.nand$1_0.Z 0.07835f
C252 v_ref vspike 0.2195f
C253 v_ref a_3544_2068# 0.137f
C254 vin ota_1stage$2_0.vp 0
C255 vin a_6854_3116# 0.21271f
C256 a_9352_5200# vdd 0.2791f
C257 vdd a_7562_3851# 1.2793f
C258 v_ref a_2248_2068# 0.01335f
C259 vmem v_th 0.01055f
C260 a_1078_602# phaseUpulse_0.monostable_0.not$1_0.in 0.00381f
C261 vin a_6164_1900# 0.21486f
C262 vdd vspike 0.90157f
C263 vdd a_3544_2068# 0.27055f
C264 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_1 0.04237f
C265 ota_1stage$2_0.vout phaseUpulse_0.conmutator_0.out 0.00815f
C266 vin a_8190_3623# 0.00184f
C267 a_n1388_602# phaseUpulse_0.vneg 0.00381f
C268 vdd a_2248_2068# 0.27536f
C269 phaseUpulse_0.vrefrac a_952_2068# 0.01389f
C270 vdd phaseUpulse_0.conmutator_0.out 0.74727f
C271 vin a_7562_3851# 0.11121f
C272 phaseUpulse_0.monostable_0.not$1_1.in v_th 0.1654f
C273 phaseUpulse_0.vrefrac phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.18679f
C274 a_n1388_602# phaseUpulse_0.monostable_0.nand$1_1.Z 0.04857f
C275 vin vspike 0.18648f
C276 phaseUpulse_0.monostable_0.nand$1_0.Z vdd 0.37216f
C277 v_ref a_8075_6021# 0.06851f
C278 a_2266_4884# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.03377f
C279 a_952_2068# vspike 0.55963f
C280 a_3544_1172# phaseUpulse_0.phi_2 0.01051f
C281 vdd a_8075_6021# 0.27918f
C282 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in 0.42262f
C283 phaseUpulse_0.phi_1 phaseUpulse_0.phi_2 0.4489f
C284 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vspike 0.04355f
C285 a_952_2068# a_2248_2068# 0.00376f
C286 a_8827_1078# vmem 0.09883f
C287 a_952_2068# phaseUpulse_0.conmutator_0.out 0.10777f
C288 a_8811_n132# vmem 0.11316f
C289 a_2583_6804# ota_1stage$2_0.vp 0.08133f
C290 a_1078_602# vdd 0.00261f
C291 a_6164_1900# a_6854_3116# 0.47928f
C292 vout phi_fire 0.57965f
C293 a_n1388_602# ota_1stage$2_0.vout 0.00427f
C294 a_2248_2068# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.00329f
C295 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.conmutator_0.out 0
C296 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.monostable_0.nand$1_1.Z 0.00251f
C297 a_n1388_602# vdd 0.00261f
C298 a_8190_3623# a_6854_3116# 0.29863f
C299 phaseUpulse_0.monostable_0.nand$1_0.Z a_952_2068# 0
C300 a_2328_3444# phaseUpulse_0.phi_2 0
C301 v_ref vmem 1.14236f
C302 phaseUpulse_0.vrefrac phaseUpulse_0.phi_int 0
C303 a_2266_4884# phaseUpulse_0.vrefrac 0.0563f
C304 a_8190_3623# a_6164_1900# 0.06628f
C305 a_7562_3851# a_6854_3116# 0.39032f
C306 conmutator$1_2.out phi_fire 0.61083f
C307 a_6854_3116# vspike 0.03458f
C308 vdd vmem 1.21265f
C309 a_7562_3851# a_6164_1900# 0.04031f
C310 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.conmutator_0.out 0.00501f
C311 phaseUpulse_0.vrefrac vspike 0.18182f
C312 a_6164_1900# vspike 0.21492f
C313 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_2 0.3513f
C314 phaseUpulse_0.vrefrac a_3544_2068# 0
C315 a_9352_5200# a_8190_3623# 0.00744f
C316 a_7562_3851# a_8190_3623# 0.17539f
C317 phaseUpulse_0.phi_1 phi_fire 0.00103f
C318 phaseUpulse_0.phi_int vspike 0.27454f
C319 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.monostable_0.not$1_3.in 0.00483f
C320 a_8190_3623# vspike 0.03541f
C321 a_3544_2068# phaseUpulse_0.phi_int 0.50615f
C322 phaseUpulse_0.vrefrac a_2248_2068# 0.10994f
C323 phaseUpulse_0.vrefrac phaseUpulse_0.conmutator_0.out 0
C324 phaseUpulse_0.monostable_0.not$1_1.in vdd 0.2269f
C325 vin vmem 0.35856f
C326 a_7562_3851# vspike 0.00374f
C327 v_th phi_fire 0.12479f
C328 a_3544_1172# phaseUpulse_0.phi_1 0.01f
C329 a_2328_3444# phi_fire 0
C330 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.phi_2 0.00112f
C331 v_rew vss 0.8189f
C332 vout vss 0.49719f
C333 vin vss 3.3876f
C334 vdd vss 92.66084f
C335 a_8811_n132# vss 0.20221f
C336 a_1078_602# vss 0.07193f
C337 a_n1388_602# vss 0.07193f
C338 conmutator$1_2.out vss 1.81382f
C339 a_3544_1172# vss 0.00446f
C340 phaseUpulse_0.monostable_0.nand$1_0.Z vss 1.12845f
C341 phaseUpulse_0.monostable_0.nand$1_1.Z vss 1.16177f
C342 a_8827_1078# vss 0.50172f
C343 phaseUpulse_0.monostable_0.not$1_1.in vss 1.45112f
C344 phaseUpulse_0.monostable_0.not$1_0.in vss 0.89571f
C345 phaseUpulse_0.monostable_0.not$1_3.in vss 1.45831f
C346 a_6854_3116# vss 1.2516f
C347 a_6164_1900# vss 2.73439f
C348 a_8190_3623# vss 2.41685f
C349 a_7562_3851# vss 0.56919f
C350 a_3544_2068# vss 0.18997f
C351 a_2248_2068# vss 0.1663f
C352 a_952_2068# vss 0.16621f
C353 vspike vss 2.59613f
C354 phaseUpulse_0.conmutator_0.out vss 0.57647f
C355 phaseUpulse_0.phi_int vss 1.53321f
C356 phaseUpulse_0.phi_2 vss 1.27584f
C357 phaseUpulse_0.phi_1 vss 1.54809f
C358 a_n872_2246# vss 0.52986f
C359 a_2328_3444# vss 1.34953f
C360 phaseUpulse_0.vneg vss 3.05036f
C361 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vss 2.76567f
C362 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn vss 1.9084f
C363 a_3790_3312# vss 1.77096f
C364 phaseUpulse_0.vrefrac vss 1.5434f
C365 a_2266_4884# vss 0.58513f
C366 a_9352_5200# vss 0.49434f
C367 v_ref vss 4.73219f
C368 phaseUpulse_0.vspike_down vss 2.28274f
C369 a_1251_5604# vss 0.93919f
C370 phaseUpulse_0.vspike_up vss 2.11982f
C371 vmem vss 4.1563f
C372 a_8075_6021# vss 0.95867f
C373 phi_fire vss 6.97034f
C374 ota_1stage$2_0.vp vss 2.52081f
C375 a_2583_6804# vss 1.42121f
C376 v_th vss 6.67973f
C377 a_4045_6672# vss 1.85283f
C378 ota_1stage$2_0.vout vss 3.78502f
C379 a_2521_8244# vss 0.71367f
C380 vmem.t0 vss 0.02433f
C381 vmem.t7 vss 0.02356f
C382 vmem.t10 vss 0.02455f
C383 vmem.n0 vss 0.02904f
C384 vmem.t4 vss 0.01517f
C385 vmem.t8 vss 0.02469f
C386 vmem.t9 vss 0.02356f
C387 vmem.n1 vss 0.04772f
C388 vmem.n2 vss 0.14288f
C389 vmem.n3 vss 0.11462f
C390 vmem.t3 vss 0.07053f
C391 vmem.t2 vss 1.1281f
C392 vmem.t11 vss 0.01984f
C393 vmem.n4 vss 0.10769f
C394 vmem.n5 vss 0.2366f
C395 vmem.t1 vss 0.02348f
C396 vmem.t5 vss 0.02444f
C397 vmem.n6 vss 0.0306f
C398 vmem.n7 vss 0.176f
C399 vmem.t6 vss 0.02348f
C400 vmem.n8 vss 0.02875f
C401 phi_fire.t9 vss 0.05802f
C402 phi_fire.t13 vss 0.05152f
C403 phi_fire.t16 vss 0.0298f
C404 phi_fire.n0 vss 0.17266f
C405 phi_fire.t6 vss 0.03827f
C406 phi_fire.n1 vss 0.10892f
C407 phi_fire.n2 vss 0.32526f
C408 phi_fire.t8 vss 0.09566f
C409 phi_fire.t11 vss 0.03827f
C410 phi_fire.n3 vss 0.37147f
C411 phi_fire.t2 vss 0.0298f
C412 phi_fire.n4 vss 0.04104f
C413 phi_fire.t15 vss 0.0357f
C414 phi_fire.n5 vss 0.19819f
C415 phi_fire.t5 vss 0.05152f
C416 phi_fire.t3 vss 0.0298f
C417 phi_fire.n6 vss 0.17266f
C418 phi_fire.t10 vss 0.03827f
C419 phi_fire.n7 vss 0.11786f
C420 phi_fire.t7 vss 0.03845f
C421 phi_fire.t12 vss 0.0298f
C422 phi_fire.n8 vss 0.03914f
C423 phi_fire.t14 vss 0.0357f
C424 phi_fire.n9 vss 0.26287f
C425 phi_fire.n10 vss 0.26273f
C426 phi_fire.t4 vss 0.05215f
C427 phi_fire.n11 vss 0.40418f
C428 phi_fire.n12 vss 1.05641f
C429 phi_fire.n13 vss 0.77893f
C430 phi_fire.t0 vss 0.06005f
C431 phi_fire.n14 vss 0.25234f
C432 phi_fire.t1 vss 0.0614f
C433 vdd.n0 vss 0.0041f
C434 vdd.n1 vss 0.01884f
C435 vdd.n2 vss 0.01025f
C436 vdd.n3 vss 0.00181f
C437 vdd.n4 vss 0.00787f
C438 vdd.n5 vss 0.00817f
C439 vdd.n6 vss 0.0067f
C440 vdd.n7 vss 0.00677f
C441 vdd.t5 vss 0.00254f
C442 vdd.n8 vss 0.00806f
C443 vdd.n9 vss 0.02142f
C444 vdd.n10 vss 0.00372f
C445 vdd.n11 vss 0.0025f
C446 vdd.n12 vss 0.01036f
C447 vdd.n13 vss 0.00669f
C448 vdd.n14 vss 0.00703f
C449 vdd.n15 vss 0.00435f
C450 vdd.n16 vss 0.00533f
C451 vdd.t4 vss 0.00254f
C452 vdd.n17 vss 0.00738f
C453 vdd.n18 vss 0.00233f
C454 vdd.n19 vss 0.00933f
C455 vdd.n20 vss 0.00977f
C456 vdd.n21 vss 0.00364f
C457 vdd.n22 vss 0.00608f
C458 vdd.n23 vss 0.00538f
C459 vdd.n24 vss 0.00372f
C460 vdd.n25 vss 0.01278f
C461 vdd.n26 vss 0.01154f
C462 vdd.t12 vss 0.03978f
C463 vdd.t13 vss 0
C464 vdd.n27 vss 0.02497f
C465 vdd.n28 vss 0.03977f
C466 vdd.n29 vss 0.02077f
C467 vdd.t38 vss 0.02416f
C468 vdd.n30 vss 0.02122f
C469 vdd.t63 vss 0.0031f
C470 vdd.t64 vss 0.02864f
C471 vdd.t62 vss 0.02928f
C472 vdd.n31 vss 0.03411f
C473 vdd.n32 vss 0.00928f
C474 vdd.n33 vss 0.05562f
C475 vdd.n34 vss 0.02629f
C476 vdd.t32 vss 0.04831f
C477 vdd.n35 vss 0.0321f
C478 vdd.t37 vss 0.0031f
C479 vdd.n36 vss 0.00236f
C480 vdd.t61 vss 0.0031f
C481 vdd.t36 vss 0.02289f
C482 vdd.t20 vss 0.02289f
C483 vdd.n37 vss 0.03406f
C484 vdd.t60 vss 0.02603f
C485 vdd.n38 vss 0.03346f
C486 vdd.n39 vss 0.01837f
C487 vdd.n40 vss 0.00715f
C488 vdd.n41 vss 0.12994f
C489 vdd.t59 vss 0.0031f
C490 vdd.n42 vss 0.00236f
C491 vdd.t57 vss 0.0031f
C492 vdd.n43 vss 0.0026f
C493 vdd.t27 vss 0.00315f
C494 vdd.t56 vss 0.03998f
C495 vdd.n44 vss 0.02271f
C496 vdd.n45 vss 0.02062f
C497 vdd.t58 vss 0.04146f
C498 vdd.t33 vss 0.03438f
C499 vdd.t40 vss 0.01935f
C500 vdd.t26 vss 0.02289f
C501 vdd.n46 vss 0.02001f
C502 vdd.n47 vss 0.02951f
C503 vdd.t35 vss 0.0031f
C504 vdd.n48 vss 0.00236f
C505 vdd.t44 vss 0.0031f
C506 vdd.n49 vss 0.0026f
C507 vdd.n50 vss 0.0398f
C508 vdd.t43 vss 0.02289f
C509 vdd.t34 vss 0.02289f
C510 vdd.n51 vss 0.03211f
C511 vdd.t25 vss 0.04189f
C512 vdd.n52 vss 0.02079f
C513 vdd.t67 vss 0.0031f
C514 vdd.n53 vss 0.0026f
C515 vdd.t29 vss 0.0031f
C516 vdd.n54 vss 0.00236f
C517 vdd.t42 vss 0.00315f
C518 vdd.t31 vss 0.00315f
C519 vdd.t66 vss 0.02306f
C520 vdd.n55 vss 0.02935f
C521 vdd.n56 vss 0.02935f
C522 vdd.t28 vss 0.03274f
C523 vdd.t41 vss 0.0292f
C524 vdd.t30 vss 0.02453f
C525 vdd.t55 vss 0.02229f
C526 vdd.n57 vss 0.02061f
C527 vdd.n58 vss 0.0353f
C528 vdd.t48 vss 0.0031f
C529 vdd.n59 vss 0.00236f
C530 vdd.t3 vss 0.0031f
C531 vdd.n60 vss 0.0026f
C532 vdd.t50 vss 0.00318f
C533 vdd.t19 vss 0.00305f
C534 vdd.n61 vss 0.00404f
C535 vdd.n62 vss 0.03401f
C536 vdd.t2 vss 0.02289f
C537 vdd.t47 vss 0.02289f
C538 vdd.n63 vss 0.03211f
C539 vdd.t18 vss 0.04207f
C540 vdd.t68 vss 0.02289f
C541 vdd.n64 vss 0.02061f
C542 vdd.t69 vss 0.0031f
C543 vdd.n65 vss 0.0026f
C544 vdd.t1 vss 0.00315f
C545 vdd.n66 vss 0.02183f
C546 vdd.t49 vss 0.03481f
C547 vdd.n67 vss 0.02726f
C548 vdd.t17 vss 0.00315f
C549 vdd.t0 vss 0.0257f
C550 vdd.t16 vss 0.02136f
C551 vdd.n68 vss 0.03966f
C552 vdd.n69 vss 0.00434f
C553 vdd.n70 vss 0.00916f
C554 vdd.n71 vss 0.00615f
C555 vdd.n72 vss 0.00391f
C556 vdd.n73 vss 0.00754f
C557 vdd.n74 vss 0.00727f
C558 vdd.n75 vss 0.0063f
C559 vdd.n76 vss 0.00637f
C560 vdd.n77 vss 0.00365f
C561 vdd.n78 vss 0.00819f
C562 vdd.n79 vss 0.00997f
C563 vdd.n80 vss 0.00266f
C564 vdd.n81 vss 0.00571f
C565 vdd.n82 vss 0.0051f
C566 vdd.n83 vss 0.00714f
C567 vdd.n84 vss 0.00554f
C568 vdd.n85 vss 0.00281f
C569 vdd.n86 vss 0.00746f
C570 vdd.n87 vss 0.00732f
C571 vdd.n88 vss 0.00443f
C572 vdd.n89 vss 0.08093f
C573 vdd.n90 vss 0.0041f
C574 vdd.n91 vss 0.01884f
C575 vdd.n92 vss 0.00538f
C576 vdd.n93 vss 0.00181f
C577 vdd.n94 vss 0.00364f
C578 vdd.n95 vss 0.00236f
C579 vdd.n96 vss 0.00608f
C580 vdd.n97 vss 0.01333f
C581 vdd.n98 vss 0.01036f
C582 vdd.n99 vss 0.0025f
C583 vdd.n100 vss 0.00787f
C584 vdd.n101 vss 0.00372f
C585 vdd.n102 vss 0.01502f
C586 vdd.n103 vss 0.02479f
C587 vdd.t54 vss 0.00457f
C588 vdd.n104 vss 0.00747f
C589 vdd.t22 vss 0.00254f
C590 vdd.n105 vss 0.00565f
C591 vdd.n106 vss 0.00736f
C592 vdd.n107 vss 0.00623f
C593 vdd.t46 vss 0.0031f
C594 vdd.t23 vss 0.11025f
C595 vdd.t21 vss 0.11025f
C596 vdd.t53 vss 0.06195f
C597 vdd.t39 vss 0.02419f
C598 vdd.n108 vss 0.02122f
C599 vdd.t65 vss 0.03003f
C600 vdd.t45 vss 0.02843f
C601 vdd.n109 vss 0.07098f
C602 vdd.n110 vss 0.03163f
C603 vdd.n111 vss 0.01071f
C604 vdd.n112 vss 0.04311f
C605 vdd.n113 vss 0.00795f
C606 vdd.n114 vss 0.00817f
C607 vdd.n115 vss 0.00792f
C608 vdd.n116 vss 0.00937f
C609 vdd.n117 vss 0.00661f
C610 vdd.n118 vss 0.0191f
C611 vdd.n119 vss 0.00915f
C612 vdd.n120 vss 0.00351f
C613 vdd.n121 vss 0.00549f
C614 vdd.n122 vss 0.00681f
C615 vdd.n123 vss 0.00817f
C616 vdd.n124 vss 0.00979f
C617 vdd.n125 vss 0.0101f
C618 vdd.t24 vss 0.00254f
C619 vdd.n126 vss 0.00743f
C620 vdd.n127 vss 0.00236f
C621 vdd.n128 vss 0.00677f
C622 vdd.n129 vss 0.0067f
C623 vdd.n130 vss 0.01025f
C624 vdd.n131 vss 0.00372f
C625 vdd.n132 vss 0.01278f
C626 vdd.n133 vss 0.01154f
C627 vdd.t15 vss 0
C628 vdd.t14 vss 0.03978f
C629 vdd.n134 vss 0.02497f
C630 vdd.n135 vss 0.03057f
C631 vdd.n136 vss 0.03588f
C632 vdd.n137 vss 0.0041f
C633 vdd.n138 vss 0.02349f
C634 vdd.n139 vss 0.01025f
C635 vdd.n140 vss 0.00181f
C636 vdd.n141 vss 0.00787f
C637 vdd.n142 vss 0.00817f
C638 vdd.n143 vss 0.0067f
C639 vdd.n144 vss 0.00677f
C640 vdd.t52 vss 0.00254f
C641 vdd.n145 vss 0.00484f
C642 vdd.t6 vss 0
C643 vdd.t7 vss 0
C644 vdd.n146 vss 0.00919f
C645 vdd.n147 vss 0.01909f
C646 vdd.n148 vss 0.01692f
C647 vdd.n149 vss 0.00372f
C648 vdd.n150 vss 0.0025f
C649 vdd.n151 vss 0.01036f
C650 vdd.n152 vss 0.00669f
C651 vdd.n153 vss 0.00703f
C652 vdd.n154 vss 0.00435f
C653 vdd.n155 vss 0.00533f
C654 vdd.t51 vss 0.00254f
C655 vdd.n156 vss 0.00738f
C656 vdd.n157 vss 0.00233f
C657 vdd.n158 vss 0.00933f
C658 vdd.n159 vss 0.00977f
C659 vdd.n160 vss 0.00364f
C660 vdd.n161 vss 0.00608f
C661 vdd.n162 vss 0.00538f
C662 vdd.n163 vss 0.00372f
C663 vdd.n164 vss 0.01692f
C664 vdd.n165 vss 0.01479f
C665 vdd.t8 vss 0
C666 vdd.t9 vss 0.00149f
C667 vdd.n166 vss 0.00942f
C668 vdd.n167 vss 0.00797f
C669 vdd.t10 vss 0.03978f
C670 vdd.t11 vss 0
C671 vdd.n168 vss 0.02497f
C672 vdd.n169 vss 0.03873f
C673 vdd.n170 vss 0.02011f
.ends

