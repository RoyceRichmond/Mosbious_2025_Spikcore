** sch_path: /foss/designs/Mosbious_2025_spiking4all/designs/libs/core_LIF_ring/LIF.sch
.subckt LIF_ring vdd vlk vout vfb vss
*.PININFO vdd:B vss:B vout:B vfb:B vlk:B
XM2 inv1 vlk vdd vdd pfet_03v3 L=50u W=0.45u nf=1 m=1
XM4 net2 inv1 vdd vdd pfet_03v3 L=0.28u W=0.45u nf=1 m=1
XM1 net1 vfb vss vss nfet_03v3 L=10u W=3u nf=1 m=1
XM3 net3 inv1 vss vss nfet_03v3 L=0.28u W=0.45u nf=1 m=1
XM5 net4 net3 vdd vdd pfet_03v3 L=0.28u W=0.45u nf=1 m=1
XM6 vout net3 vss vss nfet_03v3 L=0.28u W=0.45u nf=1 m=1
XC2 inv1 vss cap_mim_2f0fF c_width=1e-6 c_length=1e-6 m=130
.ends
