* NGSPICE file created from LIF_comp.ext - technology: gf180mcuD

.subckt LIF_comp_pex vdd vss vin v_rew vout
X0 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vss.t2 vss.t1 nfet_03v3 ad=9.15p pd=31.22u as=9.15p ps=31.22u w=15u l=0.28u
X1 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vrefrac vss.t10 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X2 a_n1388_602# ota_1stage$2_0.vout vss.t15 vss.t14 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X3 vspike a_3544_2068# v_ref vdd.t50 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X4 a_1251_6917# phaseUpulse_0.vspike_up phaseUpulse_0.vspike_up vss.t8 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X5 vss.t31 v_rew.t0 a_n872_2246# vss.t30 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X6 vspike a_2248_2068# phaseUpulse_0.vrefrac vdd.t51 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X7 vss.t29 a_4045_8037# a_2583_8169# vss.t27 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X8 a_3790_4625# a_3790_4625# vss.t39 vss.t37 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X9 a_2583_8169# v_th ota_1stage$2_0.vout vss.t85 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X10 vss.t77 v_ref v_ref vss.t76 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X11 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.not$1_3.in vdd.t2 vdd.t1 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X12 vdd.t33 vdd.t32 a_6164_1900# vss.t63 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X13 phaseUpulse_0.phi_2 phaseUpulse_0.monostable_0.not$1_0.in vdd.t57 vdd.t56 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X14 vdd.t55 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.nand$1_0.Z vdd.t54 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X15 vss.t62 phaseUpulse_0.phi_2 a_2248_2068# vss.t61 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X16 vin.t0 a_8811_n132# vmem.t1 vdd.t0 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X17 vss.t47 phi_fire.t2 a_8827_1078# vss.t46 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X18 vss.t26 phaseUpulse_0.phi_1 a_952_2068# vss.t25 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X19 v_ref a_8827_1078# conmutator$1_2.out vdd.t44 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X20 vdd.t19 v_rew.t1 a_n872_2246# vdd.t18 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X21 vdd.t31 a_2266_6197# phaseUpulse_0.vrefrac vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X22 a_4045_8037# a_4045_8037# vss.t28 vss.t27 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X23 phaseUpulse_0.phi_1 phaseUpulse_0.vneg vdd.t24 vdd.t23 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X24 v_ref a_9352_5200# vout.t1 vss.t32 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X25 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_1 vdd.t17 vdd.t16 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X26 a_7562_3851# a_7562_3851# vdd.t65 vdd.t64 pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X27 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.monostable_0.not$1_1.in cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
X28 conmutator$1_2.out phi_fire.t3 vmem.t5 vdd.t0 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X29 vdd.t22 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.nand$1_1.Z vdd.t21 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X30 vmem.t11 v_th vin.t2 vss.t84 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X31 a_8190_3623# vmem.t9 cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
X32 v_ref phi_fire.t4 conmutator$1_2.out vss.t48 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X33 vdd.t49 phaseUpulse_0.phi_2 a_2248_2068# vdd.t48 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X34 vss.t73 phaseUpulse_0.phi_int a_3544_2068# vss.t72 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X35 vdd.t43 a_2521_9609# ota_1stage$2_0.vout vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X36 a_9352_5200# phi_fire.t5 vdd.t7 vdd.t6 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X37 vin.t3 conmutator$1_2.out cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
X38 vspike phaseUpulse_0.phi_1 phaseUpulse_0.conmutator_0.out vss.t24 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X39 vmem.t10 a_8190_3623# vdd.t46 vdd.t45 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
X40 vdd.t39 vdd.t38 a_3790_4625# vss.t56 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X41 vdd.t15 phaseUpulse_0.phi_1 a_952_2068# vdd.t14 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X42 phaseUpulse_0.conmutator_0.out v_rew.t2 phaseUpulse_0.vspike_up vdd.t52 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X43 vss.t83 v_th phaseUpulse_0.monostable_0.not$1_3.in vss.t82 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
X44 phaseUpulse_0.monostable_0.nand$1_1.Z ota_1stage$2_0.vout vdd.t4 vdd.t3 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X45 conmutator$1_0.out a_8075_5978# vmem.t2 vss.t17 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X46 conmutator$1_2.out a_8827_1078# vmem.t8 vss.t57 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X47 vdd.t37 vdd.t36 a_4045_8037# vss.t68 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
X48 vdd.t9 phi_fire.t6 a_8811_n132# vdd.t8 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X49 phaseUpulse_0.phi_int phaseUpulse_0.phi_1 vss.t23 vss.t22 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X50 phaseUpulse_0.vneg phaseUpulse_0.monostable_0.not$1_3.in vss.t12 vss.t11 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X51 vspike phaseUpulse_0.phi_int v_ref vss.t71 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X52 vss.t81 v_th phaseUpulse_0.monostable_0.not$1_1.in vss.t80 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
X53 a_7562_3851# vin.t4 a_6854_3116# vss.t54 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X54 a_2328_4757# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vrefrac vss.t9 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X55 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.vneg phaseUpulse_0.vneg vss.t36 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=13u
X56 vss.t79 v_th v_th vss.t78 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.8u
X57 vspike phaseUpulse_0.phi_2 phaseUpulse_0.vrefrac vss.t9 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X58 vdd.t61 phaseUpulse_0.phi_int a_3544_2068# vdd.t60 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X59 phaseUpulse_0.phi_1 phaseUpulse_0.vneg vss.t35 vss.t34 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X60 v_ref vdd.t40 vdd.t41 vss.t55 nfet_03v3 ad=0.3355p pd=2.32u as=0.3355p ps=2.32u w=0.55u l=0.28u
X61 a_6854_3116# a_6164_1900# vss.t7 vss.t3 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X62 phaseUpulse_0.conmutator_0.out a_n872_2246# phaseUpulse_0.vspike_up vss.t86 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X63 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.monostable_0.not$1_3.in cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
X64 v_ref phi_fire.t7 vout.t3 vdd.t10 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X65 phi_fire.t1 phaseUpulse_0.phi_int vdd.t59 vdd.t58 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X66 a_1078_602# phaseUpulse_0.phi_1 vss.t21 vss.t20 nfet_03v3 ad=0.4p pd=1.8u as=0.61p ps=3.22u w=1u l=0.28u
X67 vdd.t30 a_2266_6197# a_2266_6197# vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X68 vmem.t0 a_6164_1900# vss.t6 vss.t5 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X69 vdd.t28 phi_fire.t8 a_8827_1078# vdd.t27 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X70 vdd.t63 a_7562_3851# a_8190_3623# vdd.t62 pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X71 phaseUpulse_0.phi_int phaseUpulse_0.phi_2 a_3544_1172# vdd.t47 pfet_03v3 ad=0.65p pd=3.3u as=0.42p ps=1.84u w=1u l=0.28u
X72 conmutator$1_0.out phi_fire.t9 vmem.t4 vdd.t29 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X73 a_6854_3116# vspike a_8190_3623# vss.t58 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X74 vss.t4 a_6164_1900# a_6164_1900# vss.t3 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X75 phaseUpulse_0.vspike_down a_1251_6917# a_1251_6917# vss.t19 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X76 a_2583_8169# conmutator$1_0.out a_2521_9609# vss.t18 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X77 vss.t45 phi_fire.t10 conmutator$1_0.out vss.t44 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X78 vdd.t42 a_2521_9609# a_2521_9609# vdd pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
X79 vss.t50 phi_fire.t11 a_8811_n132# vss.t49 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X80 vdd.t53 v_rew.t3 phaseUpulse_0.conmutator_0.out vss.t64 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X81 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in vdd.t67 vdd.t66 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X82 a_3544_1172# phaseUpulse_0.phi_1 vdd.t13 vdd.t12 pfet_03v3 ad=0.42p pd=1.84u as=0.65p ps=3.3u w=1u l=0.28u
X83 vout.t2 phi_fire.t12 vmem.t6 vss.t51 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X84 v_th phaseUpulse_0.vspike_down phaseUpulse_0.vspike_down vss.t13 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X85 vin.t1 phi_fire.t13 vmem.t7 vss.t52 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X86 phi_fire.t0 phaseUpulse_0.phi_int vss.t70 vss.t69 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X87 vdd.t69 a_n872_2246# phaseUpulse_0.conmutator_0.out vdd.t68 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X88 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vneg a_n1388_602# vss.t33 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X89 phaseUpulse_0.vspike_up vdd.t34 vdd.t35 vss.t53 nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
X90 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.monostable_0.not$1_0.in a_1078_602# vss.t67 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X91 vdd.t26 phi_fire.t14 a_8075_5978# vdd.t25 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X92 vspike a_952_2068# phaseUpulse_0.conmutator_0.out vdd.t5 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X93 vout.t0 a_9352_5200# vmem.t3 vdd.t20 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
X94 a_9352_5200# phi_fire.t15 vss.t41 vss.t40 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X95 a_2328_4757# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp a_2266_6197# vss.t0 nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
X96 vss.t60 phaseUpulse_0.phi_2 phaseUpulse_0.phi_int vss.t59 nfet_03v3 ad=0.61p pd=3.22u as=0.4p ps=1.8u w=1u l=0.28u
X97 vss.t43 phi_fire.t16 a_8075_5978# vss.t42 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X98 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vspike_down phaseUpulse_0.vspike_down vss.t10 nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
X99 vss.t38 a_3790_4625# a_2328_4757# vss.t37 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
X100 phaseUpulse_0.phi_2 phaseUpulse_0.monostable_0.not$1_0.in vss.t66 vss.t65 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X101 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in vss.t75 vss.t74 nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
X102 vss.t16 a_8075_5978# conmutator$1_0.out vdd.t11 pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
R0 vss.n1201 vss.n212 52569.5
R1 vss.n1200 vss.n1199 12732.4
R2 vss.n1387 vss.n442 7073.53
R3 vss.n1628 vss.n139 6997.06
R4 vss.n1117 vss.n81 6933.33
R5 vss.n212 vss.n139 6767.65
R6 vss.n734 vss.n681 6102.12
R7 vss.n799 vss.n797 4445.99
R8 vss.n1405 vss.t71 3976.47
R9 vss.t55 vss.n1117 3683.33
R10 vss.t1 vss.n401 3619.61
R11 vss.n1372 vss.t36 3441.18
R12 vss.n797 vss.n733 3319.89
R13 vss.n1105 vss.n81 3135.29
R14 vss.t1 vss.n400 2931.37
R15 vss.n733 vss.n682 2746.31
R16 vss.n1199 vss.t55 2740.2
R17 vss.n1405 vss.t36 2498.04
R18 vss.n1332 vss.n1331 2281.37
R19 vss.n1330 vss.n446 2281.37
R20 vss.n1357 vss.n442 2281.37
R21 vss.n1201 vss.n1200 2166.67
R22 vss.t69 vss.n922 2021.95
R23 vss.n1620 vss.n1619 1853.24
R24 vss.n1628 vss.n1627 1848.04
R25 vss.n1372 vss.n401 1835.29
R26 vss.n1331 vss.n1330 1822.55
R27 vss.n801 vss.n681 1429.64
R28 vss.n802 vss.n680 1314.21
R29 vss.n1094 vss.n1079 1305.17
R30 vss.n1627 vss.n140 1300
R31 vss.n1619 vss.n140 1300
R32 vss.n1095 vss.n1094 1300
R33 vss.n1096 vss.n1095 1300
R34 vss.n1096 vss.n1074 1300
R35 vss.n1104 vss.n1074 1300
R36 vss.n1105 vss.n1104 1300
R37 vss.n1333 vss.n457 1300
R38 vss.n1333 vss.n1332 1300
R39 vss.n1356 vss.n446 1300
R40 vss.n1357 vss.n1356 1300
R41 vss.t52 vss.t49 1200
R42 vss.n769 vss.n762 910.816
R43 vss.n770 vss.n769 905.739
R44 vss.n786 vss.n770 905.739
R45 vss.n786 vss.n785 905.739
R46 vss.n785 vss.n784 905.739
R47 vss.n784 vss.n771 905.739
R48 vss.n771 vss.n680 905.739
R49 vss.t40 vss.t51 862.323
R50 vss.t63 vss.n555 861.788
R51 vss.n797 vss.n796 851.777
R52 vss.t44 vss.t42 823.909
R53 vss.t49 vss.n799 781.25
R54 vss.n800 vss.t52 781.25
R55 vss.n1288 vss.n468 777
R56 vss.t59 vss.n923 740.376
R57 vss.n1017 vss.t67 740.376
R58 vss.n999 vss.t33 740.376
R59 vss.n1387 vss.n400 688.236
R60 vss.n801 vss.n800 665.625
R61 vss.n943 vss.n924 625.567
R62 vss.n979 vss.n960 625.567
R63 vss.n512 vss.n468 610.4
R64 vss.n688 vss.n687 591.159
R65 vss.n683 vss.t32 549.77
R66 vss.t17 vss.n689 498.435
R67 vss.n732 vss.t32 467.491
R68 vss.t51 vss.n683 467.491
R69 vss.t1 vss.n212 429.981
R70 vss.n689 vss.t44 423.839
R71 vss.n690 vss.t17 423.839
R72 vss.n744 vss.t46 386.286
R73 vss.n996 vss.t14 378.729
R74 vss.n923 vss.t69 367.981
R75 vss.n924 vss.t22 367.981
R76 vss.n1018 vss.t74 367.981
R77 vss.t74 vss.n1017 367.981
R78 vss.n960 vss.t20 367.981
R79 vss.n1000 vss.t11 367.981
R80 vss.t11 vss.n999 367.981
R81 vss.n690 vss.n682 361.111
R82 vss.n555 vss.n5 336.683
R83 vss.t22 vss.t59 317.935
R84 vss.t20 vss.t67 317.935
R85 vss.t14 vss.t33 317.935
R86 vss.n792 vss.n737 290.378
R87 vss.n796 vss.t46 236.606
R88 vss.n1201 vss.t36 228.376
R89 vss.n1019 vss.n1018 195.766
R90 vss.n1001 vss.n1000 195.766
R91 vss.n754 vss.t48 186.673
R92 vss.n802 vss.n801 177.596
R93 vss.n139 vss.n138 167.925
R94 vss.n754 vss.t5 162.739
R95 vss.t64 vss.t30 155.767
R96 vss.t57 vss.n681 154.762
R97 vss.n1288 vss.n1287 153.263
R98 vss.n1027 vss.n1026 150.137
R99 vss.n1019 vss.n931 150.137
R100 vss.n1009 vss.n1008 150.137
R101 vss.n1001 vss.n967 150.137
R102 vss.n168 vss.n100 139.507
R103 vss.n187 vss.n149 131.757
R104 vss.n1636 vss.n112 131.757
R105 vss.n827 vss.n826 131.125
R106 vss.n825 vss.n673 131.125
R107 vss.n835 vss.n545 131.125
R108 vss.n1658 vss.t18 129.173
R109 vss.n826 vss.n825 123.919
R110 vss.n910 vss.n548 120.415
R111 vss.n920 vss.n548 120.415
R112 vss.t86 vss.n305 119.26
R113 vss.n733 vss.n732 117.808
R114 vss.n1201 vss.n457 114.707
R115 vss.n793 vss.n792 113.279
R116 vss vss.t86 112.478
R117 vss.n1650 vss.t18 107.215
R118 vss.n147 vss.n92 107.215
R119 vss.n744 vss.t48 103.707
R120 vss.n943 vss.t65 103.034
R121 vss.n979 vss.t34 103.034
R122 vss.n1643 vss.n101 102.047
R123 vss.n109 vss.t85 102.047
R124 vss.t30 vss.n304 101.41
R125 vss.n305 vss.t64 101.41
R126 vss.n921 vss.n545 99.4241
R127 vss.n922 vss.n921 97.6466
R128 vss.n168 vss.n149 96.8805
R129 vss.n687 vss.t40 96.2357
R130 vss.t42 vss.n688 96.2357
R131 vss.n1643 vss.n100 95.5887
R132 vss.n1027 vss.t65 92.7315
R133 vss.n1009 vss.t34 92.7315
R134 vss.n1659 vss.n81 83.9631
R135 vss.n721 vss.n695 83.9245
R136 vss.n1026 vss.t80 75.0684
R137 vss.n1008 vss.t82 75.0684
R138 vss.n310 vss.n256 73.8273
R139 vss.n303 vss.n259 73.8273
R140 vss.n890 vss.n559 73.8273
R141 vss.n902 vss.n566 73.8273
R142 vss.n611 vss.n610 73.8273
R143 vss.n1688 vss.n5 73.8273
R144 vss.n827 vss.t58 73.4875
R145 vss.n673 vss.t54 73.4875
R146 vss.n835 vss.t54 73.4875
R147 vss.n1420 vss.n410 69.8337
R148 vss.n1451 vss.n1450 69.8337
R149 vss.n1478 vss.n368 69.8337
R150 vss.n1472 vss.n1471 69.8337
R151 vss.n336 vss.n328 69.8337
R152 vss.n1614 vss.n1613 69.8337
R153 vss.t78 vss.n147 65.8789
R154 vss.t13 vss.n1636 65.8789
R155 vss.n737 vss.t57 65.4153
R156 vss.n1461 vss.n1460 65.2394
R157 vss.n1521 vss.t9 65.2394
R158 vss.n1529 vss.n335 65.2394
R159 vss.n148 vss.t78 62.0037
R160 vss.n902 vss.n559 58.4129
R161 vss.n1231 vss.n529 57.196
R162 vss.n1484 vss.n1483 56.0508
R163 vss.n715 vss.n695 55.9499
R164 vss.n610 vss.n555 51.517
R165 vss.t80 vss.n1025 50.0458
R166 vss.t82 vss.n1007 50.0458
R167 vss.n793 vss.t5 49.4605
R168 vss.n1362 vss.n400 48.7
R169 vss.t24 vss.n247 47.4606
R170 vss.n921 vss.n920 46.0412
R171 vss.n844 vss.n625 45.4324
R172 vss.t1 vss.t36 43.8098
R173 vss.t8 vss.n247 41.3759
R174 vss.n259 vss.t53 41.3759
R175 vss.n852 vss.t3 41.3759
R176 vss.n890 vss.t3 41.3759
R177 vss.n1380 vss.n420 41.3491
R178 vss.n910 vss.n555 41.3191
R179 vss.n801 vss.t58 40.3463
R180 vss.n309 vss.t53 40.159
R181 vss.n921 vss.n546 38.9456
R182 vss.n1637 vss.t13 36.169
R183 vss.n407 vss.n405 35.836
R184 vss.t0 vss.n398 35.836
R185 vss.n611 vss.t63 35.697
R186 vss.t0 vss.n1441 33.9982
R187 vss.n1444 vss.t1 33.9982
R188 vss.n1541 vss.n330 31.2417
R189 vss.t37 vss.n427 30.4236
R190 vss.n301 vss.n261 30.0268
R191 vss.n297 vss.n260 30.0268
R192 vss.n1124 vss.n1065 30.0268
R193 vss.n1181 vss.n1126 30.0268
R194 vss.n876 vss.n620 29.7505
R195 vss.n889 vss.n622 29.7505
R196 vss.n867 vss.n619 29.7505
R197 vss.n891 vss.n618 29.7505
R198 vss.n851 vss.n628 29.7505
R199 vss.n1129 vss.n64 29.7505
R200 vss.n1673 vss.n61 29.7505
R201 vss.n1665 vss.n76 29.7505
R202 vss.n1128 vss.n65 29.7505
R203 vss.n1671 vss.n67 29.7505
R204 vss.n1308 vss.n460 29.7505
R205 vss.n1305 vss.n461 29.7505
R206 vss.n1321 vss.n462 29.7505
R207 vss.n497 vss.n496 29.7505
R208 vss.t85 vss.n101 29.7104
R209 vss.n1637 vss.n109 29.7104
R210 vss.n1688 vss.n6 29.6123
R211 vss.n1044 vss.n1043 29.3207
R212 vss.n852 vss.n625 28.3954
R213 vss.n715 vss.t84 27.9752
R214 vss.t84 vss.n546 27.9752
R215 vss.n755 vss.n741 27.1716
R216 vss.n791 vss.n739 27.1716
R217 vss.n1638 vss.n108 26.8952
R218 vss.n136 vss.n110 26.8952
R219 vss.n256 vss.t24 26.3672
R220 vss.n764 vss.n762 26.2571
R221 vss.n1687 vss.n7 26.2505
R222 vss.n1683 vss.n8 26.2505
R223 vss.n1148 vss.n4 26.2505
R224 vss.n1689 vss.n3 26.2505
R225 vss.n900 vss.n569 26.2505
R226 vss.n612 vss.n571 26.2505
R227 vss.n915 vss.n549 26.2505
R228 vss.n919 vss.n551 26.2505
R229 vss.n1511 vss.n351 26.2505
R230 vss.n1273 vss.n511 26.2505
R231 vss.n1202 vss.n1201 25.9616
R232 vss.n283 vss.t25 25.5559
R233 vss.n1025 vss.n931 25.0231
R234 vss.n1007 vss.n967 25.0231
R235 vss.n402 vss.n393 24.8097
R236 vss.n330 vss.n209 24.8097
R237 vss.n1650 vss.n92 24.5434
R238 vss.n775 vss.n736 24.1237
R239 vss.n710 vss.n709 23.9479
R240 vss.n706 vss.n702 23.9479
R241 vss.n720 vss.n696 23.9479
R242 vss.n723 vss.n693 23.9479
R243 vss.n1582 vss.n241 23.9479
R244 vss.n1576 vss.n238 23.9479
R245 vss.n1553 vss.n321 23.9479
R246 vss.n223 vss.n219 23.9334
R247 vss.t56 vss.n56 23.9334
R248 vss.n1380 vss.n1362 23.8908
R249 vss.n1421 vss.n1420 23.8908
R250 vss.n1435 vss.n410 23.8908
R251 vss.n1441 vss.n405 23.8908
R252 vss.n1444 vss.n398 23.8908
R253 vss.n1450 vss.n393 23.8908
R254 vss.n1451 vss.n357 23.8908
R255 vss.n1471 vss.n1461 23.8908
R256 vss.n1521 vss.n349 23.8908
R257 vss.n1529 vss.n344 23.8908
R258 vss.n1535 vss.n336 23.8908
R259 vss.n1542 vss.n328 23.8908
R260 vss.n1614 vss.n209 23.8908
R261 vss.n317 vss.n239 23.406
R262 vss.n1435 vss.t36 22.9719
R263 vss.n1035 vss.n542 22.1935
R264 vss.n1002 vss.n970 22.0137
R265 vss.n988 vss.n971 22.0137
R266 vss.n981 vss.n965 22.0137
R267 vss.n1010 vss.n963 22.0137
R268 vss.n1020 vss.n934 22.0137
R269 vss.n952 vss.n935 22.0137
R270 vss.n945 vss.n929 22.0137
R271 vss.n1028 vss.n927 22.0137
R272 vss.n1584 vss.n233 21.9051
R273 vss.n1220 vss.t76 21.9051
R274 vss.n1551 vss.n1549 21.4687
R275 vss.n477 vss.t27 21.0939
R276 vss.n721 vss.n682 20.8444
R277 vss.n1566 vss.n1563 20.7984
R278 vss.n753 vss.n742 20.0599
R279 vss.n704 vss.n0 19.7904
R280 vss.n1203 vss.n1109 19.711
R281 vss.n1616 vss.t19 19.4713
R282 vss.n1179 vss.n510 18.66
R283 vss.n1692 vss.n1691 18.4568
R284 vss.n1035 vss 18.2874
R285 vss.n1037 vss.n1036 18.0005
R286 vss.n1483 vss.t61 17.4588
R287 vss.n426 vss.n75 17.4431
R288 vss.n803 vss.n679 17.0173
R289 vss.n194 vss.n143 16.8558
R290 vss.n178 vss.n150 16.8558
R291 vss.n291 vss.n290 16.7637
R292 vss.n290 vss.n257 16.7637
R293 vss.n254 vss.n250 16.7637
R294 vss.n311 vss.n254 16.7637
R295 vss.n284 vss.n282 16.6716
R296 vss.n844 vss.n547 16.6318
R297 vss.n273 vss.n272 16.5794
R298 vss.n1606 vss.n219 16.2262
R299 vss.n1591 vss.t10 16.2262
R300 vss.n1590 vss.n229 16.2262
R301 vss.n1584 vss.n1583 16.2262
R302 vss.n1191 vss.n1190 16.211
R303 vss.n1595 vss.n1594 16.2045
R304 vss.n283 vss.n244 15.8205
R305 vss.n922 vss.n544 15.7821
R306 vss.n1421 vss.n417 15.6211
R307 vss.n368 vss.n355 15.6211
R308 vss.n1041 vss.n533 15.433
R309 vss.n1282 vss.n512 15.4156
R310 vss.n1575 vss.t8 15.0092
R311 vss.n1512 vss.n1511 14.824
R312 vss.n1216 vss.n1215 14.2095
R313 vss.n195 vss.n194 14.0926
R314 vss.n202 vss.n201 14.0926
R315 vss.n1620 vss.n202 14.0926
R316 vss.n178 vss.n177 14.0926
R317 vss.n119 vss.n114 14.0926
R318 vss.n1629 vss.n119 14.0926
R319 vss.n1514 vss.n1512 14.0926
R320 vss.n1190 vss.n1189 13.8163
R321 vss.n1484 vss.n357 13.7834
R322 vss.n1542 vss.n1541 13.7834
R323 vss.n1115 vss.n84 13.7242
R324 vss.n1652 vss.n88 13.7242
R325 vss.n1285 vss.n512 13.7242
R326 vss.n282 vss.n278 13.3558
R327 vss.n1657 vss.n84 13.3558
R328 vss.n1653 vss.n1652 13.3558
R329 vss.n1652 vss.n1651 13.3558
R330 vss.n1649 vss.n84 13.3558
R331 vss.n1119 vss.t77 13.2942
R332 vss.n837 vss.n626 13.2637
R333 vss.n647 vss.n627 13.2637
R334 vss.n666 vss.n662 13.2637
R335 vss.n834 vss.n631 13.2637
R336 vss.n853 vss.n624 13.2637
R337 vss.n809 vss.n808 13.2637
R338 vss.n837 vss.n836 13.2637
R339 vss.n808 vss.n667 13.2637
R340 vss.n828 vss.n666 13.2637
R341 vss.n1087 vss.n71 13.2637
R342 vss.n1073 vss.n82 13.2637
R343 vss.n1646 vss.n1645 13.2637
R344 vss.n1073 vss.n74 13.2637
R345 vss.n1667 vss.n73 13.2637
R346 vss.n1642 vss.n102 13.2637
R347 vss.n1660 vss.n79 13.2637
R348 vss.n104 vss.n102 13.2637
R349 vss.n1645 vss.n1644 13.2637
R350 vss.n287 vss.n254 13.2637
R351 vss.n290 vss.n289 13.2637
R352 vss.n273 vss.n249 13.2637
R353 vss.n1109 vss.n1066 13.2637
R354 vss.n1190 vss.n1111 13.2637
R355 vss.n1341 vss.n452 13.2637
R356 vss.n1329 vss.n449 13.2637
R357 vss.n456 vss.n403 13.2637
R358 vss.n1443 vss.n354 13.2637
R359 vss.n354 vss.n350 13.2637
R360 vss.n1569 vss.n1561 13.2637
R361 vss.n1562 vss.n214 12.9873
R362 vss.n476 vss.n474 12.9873
R363 vss.n420 vss.n417 12.8645
R364 vss.n921 vss.n547 12.5754
R365 vss.n1672 vss.n66 12.1697
R366 vss.n525 vss.n522 11.9968
R367 vss.n536 vss.n530 11.8821
R368 vss.n1213 vss.n526 11.8821
R369 vss.n304 vss.n303 11.7641
R370 vss.n90 vss.t79 11.5442
R371 vss.n1593 vss.t19 11.3585
R372 vss.n732 vss 11.0681
R373 vss.n407 vss.t36 11.0268
R374 vss.t1 vss.n402 11.0268
R375 vss.n749 vss.t6 11.0113
R376 vss.n1233 vss.n526 10.9833
R377 vss.n1230 vss.n530 10.9833
R378 vss.n1280 vss.n1279 10.8187
R379 vss.n1316 vss.n465 10.8187
R380 vss.n1314 vss.n1313 10.8187
R381 vss.n490 vss.n486 10.8187
R382 vss.n494 vss.n492 10.8187
R383 vss.n503 vss.n482 10.8187
R384 vss.n1293 vss.n1292 10.8187
R385 vss.n1561 vss.n318 10.7963
R386 vss.n282 vss.n281 10.5926
R387 vss.n731 vss.n683 10.59
R388 vss.n726 vss.n690 10.59
R389 vss.n727 vss.n689 10.59
R390 vss.n1013 vss.n960 10.59
R391 vss.n1031 vss.n924 10.59
R392 vss.n1541 vss.n1540 10.59
R393 vss.n306 vss.n305 10.59
R394 vss.n309 vss.n308 10.59
R395 vss.n1410 vss.n420 10.59
R396 vss.n794 vss.n793 10.59
R397 vss.n800 vss.n542 10.59
R398 vss.n1575 vss.n244 10.5472
R399 vss.n1220 vss.n1063 10.5472
R400 vss.n478 vss.n477 10.5472
R401 vss.n1399 vss.n427 10.5472
R402 vss.n1393 vss.n435 10.5472
R403 vss.n525 vss.n507 10.5005
R404 vss.n646 vss.n645 10.4483
R405 vss.n1093 vss.n1080 10.4483
R406 vss.n1343 vss.n1342 10.4483
R407 vss.n1599 vss.n1598 10.4136
R408 vss.n1226 vss.n533 10.4084
R409 vss.n687 vss.n684 10.4005
R410 vss.n688 vss.n685 10.4005
R411 vss.n923 vss.n543 10.4005
R412 vss.n1025 vss.n1024 10.4005
R413 vss.n1017 vss.n1016 10.4005
R414 vss.n1007 vss.n1006 10.4005
R415 vss.n999 vss.n998 10.4005
R416 vss.n304 vss.n258 10.4005
R417 vss.n1411 vss.n402 10.4005
R418 vss.n1056 vss.n1055 10.4005
R419 vss.n796 vss.n795 10.4005
R420 vss.n799 vss.n798 10.4005
R421 vss.n1583 vss.t25 10.1415
R422 vss.n1212 vss.n1211 10.1415
R423 vss.n1286 vss.n510 10.1415
R424 vss.n1544 vss.n325 10.1321
R425 vss.n1574 vss.n317 10.0201
R426 vss.n1574 vss.n318 9.94896
R427 vss.n1626 vss.n119 9.85576
R428 vss.n202 vss.n141 9.85576
R429 vss.n180 vss.n178 9.85576
R430 vss.n194 vss.n193 9.85576
R431 vss.n1512 vss.n1509 9.85576
R432 vss.n1672 vss.n63 9.7359
R433 vss.n1303 vss.t27 9.7359
R434 vss.n72 vss.t28 9.54445
R435 vss.n450 vss.t39 9.54445
R436 vss.n658 vss.t4 9.54445
R437 vss.n1675 vss.t29 9.54326
R438 vss.n1319 vss.t38 9.54326
R439 vss.n893 vss.t7 9.54326
R440 vss.n1687 vss.n8 9.39524
R441 vss.n1681 vss.n1680 9.39524
R442 vss.n1678 vss.n58 9.39524
R443 vss.n1136 vss.n1135 9.39524
R444 vss.n1174 vss.n1173 9.39524
R445 vss.n1171 vss.n1168 9.39524
R446 vss.n1166 vss.n1139 9.39524
R447 vss.n1161 vss.n1160 9.39524
R448 vss.n1158 vss.n1144 9.39524
R449 vss.n1151 vss.n1150 9.39524
R450 vss.n1689 vss.n4 9.39524
R451 vss.n52 vss.n50 9.39524
R452 vss.n50 vss.n49 9.39524
R453 vss.n46 vss.n45 9.39524
R454 vss.n43 vss.n12 9.39524
R455 vss.n39 vss.n37 9.39524
R456 vss.n35 vss.n14 9.39524
R457 vss.n31 vss.n29 9.39524
R458 vss.n27 vss.n16 9.39524
R459 vss.n23 vss.n21 9.39524
R460 vss.n19 vss.n3 9.39524
R461 vss.n709 vss.n708 9.39524
R462 vss.n716 vss.n696 9.39524
R463 vss.n716 vss.n698 9.39524
R464 vss.n702 vss.n698 9.39524
R465 vss.n720 vss.n694 9.39524
R466 vss.n714 vss.n693 9.39524
R467 vss.n714 vss.n699 9.39524
R468 vss.n710 vss.n699 9.39524
R469 vss.n612 vss.n569 9.39524
R470 vss.n588 vss.n571 9.39524
R471 vss.n608 vss.n589 9.39524
R472 vss.n604 vss.n603 9.39524
R473 vss.n600 vss.n599 9.39524
R474 vss.n596 vss.n595 9.39524
R475 vss.n592 vss.n591 9.39524
R476 vss.n582 vss.n574 9.39524
R477 vss.n578 vss.n577 9.39524
R478 vss.n911 vss.n554 9.39524
R479 vss.n912 vss.n911 9.39524
R480 vss.n912 vss.n549 9.39524
R481 vss.n568 vss.n567 9.39524
R482 vss.n895 vss.n567 9.39524
R483 vss.n858 vss.n857 9.39524
R484 vss.n862 vss.n861 9.39524
R485 vss.n871 vss.n870 9.39524
R486 vss.n885 vss.n884 9.39524
R487 vss.n882 vss.n881 9.39524
R488 vss.n904 vss.n558 9.39524
R489 vss.n909 vss.n556 9.39524
R490 vss.n909 vss.n550 9.39524
R491 vss.n919 vss.n550 9.39524
R492 vss.n992 vss.n991 9.39524
R493 vss.n966 vss.n965 9.39524
R494 vss.n985 vss.n966 9.39524
R495 vss.n985 vss.n971 9.39524
R496 vss.n977 vss.n975 9.39524
R497 vss.n1010 vss.n964 9.39524
R498 vss.n1003 vss.n964 9.39524
R499 vss.n1003 vss.n1002 9.39524
R500 vss.n956 vss.n955 9.39524
R501 vss.n930 vss.n929 9.39524
R502 vss.n949 vss.n930 9.39524
R503 vss.n949 vss.n935 9.39524
R504 vss.n941 vss.n939 9.39524
R505 vss.n1028 vss.n928 9.39524
R506 vss.n1021 vss.n928 9.39524
R507 vss.n1021 vss.n1020 9.39524
R508 vss.n655 vss.n626 9.39524
R509 vss.n655 vss.n620 9.39524
R510 vss.n878 vss.n622 9.39524
R511 vss.n627 vss.n621 9.39524
R512 vss.n889 vss.n621 9.39524
R513 vss.n833 vss.n662 9.39524
R514 vss.n834 vss.n833 9.39524
R515 vss.n854 vss.n853 9.39524
R516 vss.n854 vss.n619 9.39524
R517 vss.n865 vss.n618 9.39524
R518 vss.n851 vss.n617 9.39524
R519 vss.n891 vss.n617 9.39524
R520 vss.n809 vss.n660 9.39524
R521 vss.n836 vss.n660 9.39524
R522 vss.n804 vss.n803 9.39524
R523 vss.n804 vss.n667 9.39524
R524 vss.n764 vss.n665 9.39524
R525 vss.n828 vss.n665 9.39524
R526 vss.n768 vss.n763 9.39524
R527 vss.n768 vss.n760 9.39524
R528 vss.n787 vss.n760 9.39524
R529 vss.n755 vss.n738 9.39524
R530 vss.n791 vss.n738 9.39524
R531 vss.n746 vss.n742 9.39524
R532 vss.n70 vss.n64 9.39524
R533 vss.n71 vss.n70 9.39524
R534 vss.n1177 vss.n1129 9.39524
R535 vss.n1673 vss.n62 9.39524
R536 vss.n1665 vss.n62 9.39524
R537 vss.n96 vss.n82 9.39524
R538 vss.n1646 vss.n96 9.39524
R539 vss.n1153 vss.n65 9.39524
R540 vss.n1140 vss.n1128 9.39524
R541 vss.n1671 vss.n68 9.39524
R542 vss.n1667 vss.n68 9.39524
R543 vss.n1642 vss.n103 9.39524
R544 vss.n1638 vss.n103 9.39524
R545 vss.n1660 vss.n80 9.39524
R546 vss.n104 vss.n80 9.39524
R547 vss.n1644 vss.n98 9.39524
R548 vss.n110 vss.n98 9.39524
R549 vss.n127 vss.n126 9.39524
R550 vss.n131 vss.n130 9.39524
R551 vss.n135 vss.n124 9.39524
R552 vss.n284 vss.n248 9.39524
R553 vss.n291 vss.n248 9.39524
R554 vss.n296 vss.n257 9.39524
R555 vss.n297 vss.n296 9.39524
R556 vss.n316 vss.n249 9.39524
R557 vss.n316 vss.n250 9.39524
R558 vss.n311 vss.n255 9.39524
R559 vss.n261 vss.n255 9.39524
R560 vss.n275 vss.n274 9.39524
R561 vss.n1203 vss.n1110 9.39524
R562 vss.n1209 vss.n1065 9.39524
R563 vss.n1209 vss.n1066 9.39524
R564 vss.n1181 vss.n1064 9.39524
R565 vss.n1191 vss.n1064 9.39524
R566 vss.n1187 vss.n1184 9.39524
R567 vss.n1197 vss.n1111 9.39524
R568 vss.n1657 vss.n85 9.39524
R569 vss.n1626 vss.n1625 9.39524
R570 vss.n1625 vss.n141 9.39524
R571 vss.n1651 vss.n89 9.39524
R572 vss.n188 vss.n89 9.39524
R573 vss.n188 vss.n143 9.39524
R574 vss.n196 vss.n195 9.39524
R575 vss.n196 vss.n111 9.39524
R576 vss.n201 vss.n111 9.39524
R577 vss.n1620 vss.n1618 9.39524
R578 vss.n1618 vss.n203 9.39524
R579 vss.n281 vss.n203 9.39524
R580 vss.n180 vss.n179 9.39524
R581 vss.n1649 vss.n93 9.39524
R582 vss.n186 vss.n93 9.39524
R583 vss.n186 vss.n150 9.39524
R584 vss.n177 vss.n113 9.39524
R585 vss.n1635 vss.n113 9.39524
R586 vss.n1635 vss.n114 9.39524
R587 vss.n1629 vss.n120 9.39524
R588 vss.n267 vss.n120 9.39524
R589 vss.n272 vss.n267 9.39524
R590 vss.n1226 vss.n1225 9.39524
R591 vss.n1225 vss.n534 9.39524
R592 vss.n1053 vss.n534 9.39524
R593 vss.n1053 vss.n1047 9.39524
R594 vss.n1047 vss.n428 9.39524
R595 vss.n1398 vss.n428 9.39524
R596 vss.n1398 vss.n429 9.39524
R597 vss.n1371 vss.n429 9.39524
R598 vss.n1371 vss.n1367 9.39524
R599 vss.n1374 vss.n414 9.39524
R600 vss.n1422 vss.n414 9.39524
R601 vss.n1423 vss.n1422 9.39524
R602 vss.n1431 vss.n1423 9.39524
R603 vss.n1431 vss.n1430 9.39524
R604 vss.n1430 vss.n1424 9.39524
R605 vss.n1424 vss.n362 9.39524
R606 vss.n1482 vss.n362 9.39524
R607 vss.n1482 vss.n363 9.39524
R608 vss.n1470 vss.n363 9.39524
R609 vss.n1470 vss.n1462 9.39524
R610 vss.n1462 vss.n337 9.39524
R611 vss.n1534 vss.n337 9.39524
R612 vss.n1534 vss.n338 9.39524
R613 vss.n338 vss.n213 9.39524
R614 vss.n1612 vss.n213 9.39524
R615 vss.n1612 vss.n214 9.39524
R616 vss.n1222 vss.n536 9.39524
R617 vss.n1222 vss.n1221 9.39524
R618 vss.n1221 vss.n537 9.39524
R619 vss.n537 vss.n475 9.39524
R620 vss.n475 vss.n432 9.39524
R621 vss.n1395 vss.n432 9.39524
R622 vss.n1395 vss.n1394 9.39524
R623 vss.n1394 vss.n433 9.39524
R624 vss.n1365 vss.n433 9.39524
R625 vss.n1379 vss.n1363 9.39524
R626 vss.n1379 vss.n411 9.39524
R627 vss.n1434 vss.n411 9.39524
R628 vss.n1434 vss.n406 9.39524
R629 vss.n406 vss.n399 9.39524
R630 vss.n399 vss.n394 9.39524
R631 vss.n394 vss.n366 9.39524
R632 vss.n1479 vss.n366 9.39524
R633 vss.n1479 vss.n367 9.39524
R634 vss.n1467 vss.n367 9.39524
R635 vss.n1467 vss.n343 9.39524
R636 vss.n1530 vss.n343 9.39524
R637 vss.n1531 vss.n1530 9.39524
R638 vss.n1531 vss.n329 9.39524
R639 vss.n329 vss.n210 9.39524
R640 vss.n210 vss.n205 9.39524
R641 vss.n1607 vss.n205 9.39524
R642 vss.n1607 vss.n217 9.39524
R643 vss.n1214 vss.n1213 9.39524
R644 vss.n1219 vss.n1214 9.39524
R645 vss.n1551 vss.n1550 9.39524
R646 vss.n1550 vss.n320 9.39524
R647 vss.n320 vss.n239 9.39524
R648 vss.n1578 vss.n241 9.39524
R649 vss.n1554 vss.n1553 9.39524
R650 vss.n1555 vss.n1554 9.39524
R651 vss.n1555 vss.n238 9.39524
R652 vss.n1494 vss.n321 9.39524
R653 vss.n1514 vss.n1513 9.39524
R654 vss.n1513 vss.n240 9.39524
R655 vss.n1582 vss.n240 9.39524
R656 vss.n1326 vss.n460 9.39524
R657 vss.n1326 vss.n452 9.39524
R658 vss.n1305 vss.n471 9.39524
R659 vss.n1325 vss.n461 9.39524
R660 vss.n1325 vss.n462 9.39524
R661 vss.n500 vss.n474 9.39524
R662 vss.n496 vss.n458 9.39524
R663 vss.n1329 vss.n458 9.39524
R664 vss.n1442 vss.n403 9.39524
R665 vss.n1443 vss.n1442 9.39524
R666 vss.n1520 vss.n350 9.39524
R667 vss.n1520 vss.n351 9.39524
R668 vss.n1506 vss.n1497 9.39524
R669 vss.n1504 vss.n1500 9.39524
R670 vss.n1287 vss.n507 9.39524
R671 vss.n1285 vss.n511 9.39524
R672 vss.n1271 vss.n1270 9.39524
R673 vss.n1270 vss.n514 9.39524
R674 vss.n1266 vss.n1264 9.39524
R675 vss.n1262 vss.n516 9.39524
R676 vss.n1258 vss.n1256 9.39524
R677 vss.n1254 vss.n518 9.39524
R678 vss.n1250 vss.n1248 9.39524
R679 vss.n1246 vss.n520 9.39524
R680 vss.n1242 vss.n1240 9.39524
R681 vss.n1238 vss.n522 9.39524
R682 vss.n1044 vss.n539 9.39524
R683 vss.n1062 vss.n539 9.39524
R684 vss.n1062 vss.n540 9.39524
R685 vss.n1057 vss.n540 9.39524
R686 vss.n1057 vss.n425 9.39524
R687 vss.n1400 vss.n425 9.39524
R688 vss.n1400 vss.n423 9.39524
R689 vss.n1404 vss.n423 9.39524
R690 vss.n1404 vss.n422 9.39524
R691 vss.n1407 vss.n418 9.39524
R692 vss.n1419 vss.n418 9.39524
R693 vss.n1419 vss.n419 9.39524
R694 vss.n1415 vss.n419 9.39524
R695 vss.n1415 vss.n1414 9.39524
R696 vss.n1414 vss.n392 9.39524
R697 vss.n1452 vss.n392 9.39524
R698 vss.n1452 vss.n361 9.39524
R699 vss.n389 vss.n361 9.39524
R700 vss.n1459 vss.n389 9.39524
R701 vss.n1459 vss.n390 9.39524
R702 vss.n390 vss.n333 9.39524
R703 vss.n1536 vss.n333 9.39524
R704 vss.n1537 vss.n1536 9.39524
R705 vss.n1538 vss.n1537 9.39524
R706 vss.n1538 vss.n211 9.39524
R707 vss.n1594 vss.n211 9.39524
R708 vss.n1569 vss.n1568 9.39524
R709 vss.n1593 vss.n218 9.33025
R710 vss.n1055 vss.n63 9.33025
R711 vss.n478 vss.t72 9.33025
R712 vss.n526 vss.n525 9.2936
R713 vss.n533 vss.n530 9.2936
R714 vss.n962 vss.t83 9.08339
R715 vss.n926 vss.t81 9.08339
R716 vss.n996 vss.t15 9.00997
R717 vss.n1014 vss.t21 9.00997
R718 vss.n1033 vss.t60 9.00997
R719 vss.n1032 vss.t23 9.00997
R720 vss.n798 vss.t50 8.98866
R721 vss.n684 vss.t43 8.98866
R722 vss.n685 vss.t41 8.98866
R723 vss.n795 vss.t47 8.98866
R724 vss.n1411 vss.t62 8.98866
R725 vss.n258 vss.t31 8.98866
R726 vss.n1056 vss.t73 8.98866
R727 vss.n998 vss.t12 8.98025
R728 vss.n1006 vss.t35 8.98025
R729 vss.n1016 vss.t75 8.98025
R730 vss.n543 vss.t70 8.98025
R731 vss.n1024 vss.t66 8.98025
R732 vss.n1598 vss.t26 8.97572
R733 vss.n1545 vss.n206 8.94494
R734 vss.n1180 vss.n1063 8.92461
R735 vss.n472 vss.n66 8.92461
R736 vss.n686 vss.t45 8.8205
R737 vss vss.t16 8.53506
R738 vss.n1599 vss.n224 8.51897
R739 vss.n1054 vss.n466 8.51897
R740 vss.n1306 vss.n472 8.51897
R741 vss.n1472 vss.n355 8.27022
R742 vss.n1600 vss.n1599 7.70769
R743 vss.n274 vss.n273 7.36892
R744 vss.n1184 vss.n1109 7.36892
R745 vss.n1478 vss.t61 6.4325
R746 vss.n1230 vss.n527 6.15567
R747 vss.n228 vss.n217 5.9592
R748 vss.n1311 vss.n468 5.83383
R749 vss.n212 vss.n204 5.67948
R750 vss.t63 vss.n566 5.67948
R751 vss.t68 vss.n528 5.67948
R752 vss.n753 vss.n743 5.40959
R753 vss.n743 vss.n736 5.40959
R754 vss.n1040 vss.t68 5.27384
R755 vss.n509 vss.t56 5.27384
R756 vss.n1126 vss.n1120 5.22638
R757 vss.n1020 vss.n933 5.2005
R758 vss.n1020 vss.n1019 5.2005
R759 vss.n1022 vss.n1021 5.2005
R760 vss.n1021 vss.n931 5.2005
R761 vss.n932 vss.n928 5.2005
R762 vss.n1026 vss.n928 5.2005
R763 vss.n1029 vss.n1028 5.2005
R764 vss.n1028 vss.n1027 5.2005
R765 vss.n927 vss.n925 5.2005
R766 vss.n941 vss.n940 5.2005
R767 vss.n939 vss.n938 5.2005
R768 vss.n946 vss.n945 5.2005
R769 vss.n953 vss.n952 5.2005
R770 vss.n955 vss.n954 5.2005
R771 vss.n957 vss.n956 5.2005
R772 vss.n958 vss.n934 5.2005
R773 vss.n951 vss.n935 5.2005
R774 vss.n1019 vss.n935 5.2005
R775 vss.n950 vss.n949 5.2005
R776 vss.n949 vss.n931 5.2005
R777 vss.n948 vss.n930 5.2005
R778 vss.n1026 vss.n930 5.2005
R779 vss.n947 vss.n929 5.2005
R780 vss.n1027 vss.n929 5.2005
R781 vss.n1002 vss.n969 5.2005
R782 vss.n1002 vss.n1001 5.2005
R783 vss.n1004 vss.n1003 5.2005
R784 vss.n1003 vss.n967 5.2005
R785 vss.n968 vss.n964 5.2005
R786 vss.n1008 vss.n964 5.2005
R787 vss.n1011 vss.n1010 5.2005
R788 vss.n1010 vss.n1009 5.2005
R789 vss.n963 vss.n961 5.2005
R790 vss.n977 vss.n976 5.2005
R791 vss.n975 vss.n974 5.2005
R792 vss.n982 vss.n981 5.2005
R793 vss.n989 vss.n988 5.2005
R794 vss.n991 vss.n990 5.2005
R795 vss.n993 vss.n992 5.2005
R796 vss.n994 vss.n970 5.2005
R797 vss.n987 vss.n971 5.2005
R798 vss.n1001 vss.n971 5.2005
R799 vss.n986 vss.n985 5.2005
R800 vss.n985 vss.n967 5.2005
R801 vss.n984 vss.n966 5.2005
R802 vss.n1008 vss.n966 5.2005
R803 vss.n983 vss.n965 5.2005
R804 vss.n1009 vss.n965 5.2005
R805 vss.n1603 vss.n220 5.2005
R806 vss.n220 vss.n219 5.2005
R807 vss.n222 vss.n221 5.2005
R808 vss.n224 vss.n222 5.2005
R809 vss.n1587 vss.n230 5.2005
R810 vss.n230 vss.n229 5.2005
R811 vss.n232 vss.n231 5.2005
R812 vss.n1583 vss.n232 5.2005
R813 vss.n1572 vss.n246 5.2005
R814 vss.n1575 vss.n246 5.2005
R815 vss.n1574 vss.n1573 5.2005
R816 vss.n1575 vss.n1574 5.2005
R817 vss.n1559 vss.n245 5.2005
R818 vss.n1575 vss.n245 5.2005
R819 vss.n1552 vss.n1551 5.2005
R820 vss.n1551 vss.n219 5.2005
R821 vss.n1550 vss.n319 5.2005
R822 vss.n1550 vss.n224 5.2005
R823 vss.n1556 vss.n320 5.2005
R824 vss.n320 vss.n229 5.2005
R825 vss.n1557 vss.n239 5.2005
R826 vss.n1583 vss.n239 5.2005
R827 vss.n1515 vss.n1514 5.2005
R828 vss.n1514 vss.n219 5.2005
R829 vss.n1513 vss.n1492 5.2005
R830 vss.n1513 vss.n224 5.2005
R831 vss.n242 vss.n240 5.2005
R832 vss.n240 vss.n229 5.2005
R833 vss.n1582 vss.n1581 5.2005
R834 vss.n1583 vss.n1582 5.2005
R835 vss.n1509 vss.n1508 5.2005
R836 vss.n1495 vss.n1494 5.2005
R837 vss.n1502 vss.n321 5.2005
R838 vss.n321 vss.n204 5.2005
R839 vss.n1576 vss.n243 5.2005
R840 vss.n1579 vss.n1578 5.2005
R841 vss.n1580 vss.n241 5.2005
R842 vss.n1575 vss.n241 5.2005
R843 vss.n1557 vss.n238 5.2005
R844 vss.n1583 vss.n238 5.2005
R845 vss.n1556 vss.n1555 5.2005
R846 vss.n1555 vss.n229 5.2005
R847 vss.n1554 vss.n319 5.2005
R848 vss.n1554 vss.n224 5.2005
R849 vss.n1553 vss.n1552 5.2005
R850 vss.n1553 vss.n219 5.2005
R851 vss.n1549 vss.n1548 5.2005
R852 vss.n1546 vss.n204 5.2005
R853 vss.n1586 vss.n1585 5.2005
R854 vss.n1585 vss.n1584 5.2005
R855 vss.n1589 vss.n1588 5.2005
R856 vss.n1590 vss.n1589 5.2005
R857 vss.n1602 vss.n1601 5.2005
R858 vss.n1601 vss.n1600 5.2005
R859 vss.n1605 vss.n1604 5.2005
R860 vss.n1606 vss.n1605 5.2005
R861 vss.n1615 vss.n207 5.2005
R862 vss.n1616 vss.n1615 5.2005
R863 vss.n1566 vss.n1565 5.2005
R864 vss.n1568 vss.n1560 5.2005
R865 vss.n1570 vss.n1569 5.2005
R866 vss.n1569 vss.n244 5.2005
R867 vss.n1584 vss.n237 5.2005
R868 vss.n1590 vss.n228 5.2005
R869 vss.n217 vss.n216 5.2005
R870 vss.n1600 vss.n217 5.2005
R871 vss.n1608 vss.n1607 5.2005
R872 vss.n1607 vss.n1606 5.2005
R873 vss.n1610 vss.n205 5.2005
R874 vss.n1616 vss.n205 5.2005
R875 vss.n1609 vss.n214 5.2005
R876 vss.n1593 vss.n214 5.2005
R877 vss.n1596 vss.n1595 5.2005
R878 vss.n234 vss.n227 5.2005
R879 vss.n120 vss.n118 5.2005
R880 vss.n1617 vss.n120 5.2005
R881 vss.n268 vss.n267 5.2005
R882 vss.n267 vss.n218 5.2005
R883 vss.n272 vss.n271 5.2005
R884 vss.n272 vss.n223 5.2005
R885 vss.n285 vss.n284 5.2005
R886 vss.n284 vss.n283 5.2005
R887 vss.n286 vss.n248 5.2005
R888 vss.t8 vss.n248 5.2005
R889 vss.n292 vss.n291 5.2005
R890 vss.n291 vss.n247 5.2005
R891 vss.n294 vss.n257 5.2005
R892 vss.n310 vss.n257 5.2005
R893 vss.n296 vss.n295 5.2005
R894 vss.n296 vss.t53 5.2005
R895 vss.n298 vss.n297 5.2005
R896 vss.n297 vss.n259 5.2005
R897 vss.n278 vss.n277 5.2005
R898 vss.n276 vss.n275 5.2005
R899 vss.n274 vss.n266 5.2005
R900 vss.n274 vss.n233 5.2005
R901 vss.n251 vss.n249 5.2005
R902 vss.n283 vss.n249 5.2005
R903 vss.n316 vss.n315 5.2005
R904 vss.t8 vss.n316 5.2005
R905 vss.n314 vss.n250 5.2005
R906 vss.n250 vss.n247 5.2005
R907 vss.n312 vss.n311 5.2005
R908 vss.n311 vss.n310 5.2005
R909 vss.n255 vss.n253 5.2005
R910 vss.t53 vss.n255 5.2005
R911 vss.n262 vss.n261 5.2005
R912 vss.n261 vss.n259 5.2005
R913 vss.n301 vss.n300 5.2005
R914 vss.n299 vss.n260 5.2005
R915 vss.n287 vss.n252 5.2005
R916 vss.n289 vss.n263 5.2005
R917 vss.n1618 vss.n200 5.2005
R918 vss.n1618 vss.n1617 5.2005
R919 vss.n279 vss.n203 5.2005
R920 vss.n218 vss.n203 5.2005
R921 vss.n281 vss.n280 5.2005
R922 vss.n281 vss.n223 5.2005
R923 vss.n1630 vss.n1629 5.2005
R924 vss.n1629 vss.n1628 5.2005
R925 vss.n1623 vss.n141 5.2005
R926 vss.n1619 vss.n141 5.2005
R927 vss.n1625 vss.n1624 5.2005
R928 vss.n1625 vss.n140 5.2005
R929 vss.n1626 vss.n117 5.2005
R930 vss.n1627 vss.n1626 5.2005
R931 vss.n1621 vss.n1620 5.2005
R932 vss.n1649 vss.n1648 5.2005
R933 vss.n1650 vss.n1649 5.2005
R934 vss.n95 vss.n93 5.2005
R935 vss.n147 vss.n93 5.2005
R936 vss.n186 vss.n185 5.2005
R937 vss.n187 vss.n186 5.2005
R938 vss.n183 vss.n150 5.2005
R939 vss.n150 vss.n149 5.2005
R940 vss.n177 vss.n176 5.2005
R941 vss.n177 vss.n101 5.2005
R942 vss.n174 vss.n113 5.2005
R943 vss.n113 vss.n109 5.2005
R944 vss.n1635 vss.n1634 5.2005
R945 vss.n1636 vss.n1635 5.2005
R946 vss.n1633 vss.n114 5.2005
R947 vss.n114 vss.n112 5.2005
R948 vss.n1654 vss.n1653 5.2005
R949 vss.n1655 vss.n85 5.2005
R950 vss.n1657 vss.n1656 5.2005
R951 vss.n1658 vss.n1657 5.2005
R952 vss.n193 vss.n192 5.2005
R953 vss.n179 vss.n145 5.2005
R954 vss.n181 vss.n180 5.2005
R955 vss.n180 vss.n100 5.2005
R956 vss.n1651 vss.n91 5.2005
R957 vss.n1651 vss.n1650 5.2005
R958 vss.n146 vss.n89 5.2005
R959 vss.n147 vss.n89 5.2005
R960 vss.n189 vss.n188 5.2005
R961 vss.n188 vss.n187 5.2005
R962 vss.n190 vss.n143 5.2005
R963 vss.n149 vss.n143 5.2005
R964 vss.n195 vss.n142 5.2005
R965 vss.n195 vss.n101 5.2005
R966 vss.n197 vss.n196 5.2005
R967 vss.n196 vss.n109 5.2005
R968 vss.n198 vss.n111 5.2005
R969 vss.n1636 vss.n111 5.2005
R970 vss.n201 vss.n199 5.2005
R971 vss.n201 vss.n112 5.2005
R972 vss.n136 vss.n116 5.2005
R973 vss.n135 vss.n134 5.2005
R974 vss.n133 vss.n124 5.2005
R975 vss.n132 vss.n131 5.2005
R976 vss.n130 vss.n129 5.2005
R977 vss.n128 vss.n127 5.2005
R978 vss.n126 vss.n125 5.2005
R979 vss.n108 vss.n107 5.2005
R980 vss.n1661 vss.n1660 5.2005
R981 vss.n1660 vss.n1659 5.2005
R982 vss.n80 vss.n78 5.2005
R983 vss.t18 vss.n80 5.2005
R984 vss.n105 vss.n104 5.2005
R985 vss.n104 vss.n92 5.2005
R986 vss.n1642 vss.n1641 5.2005
R987 vss.n1643 vss.n1642 5.2005
R988 vss.n1640 vss.n103 5.2005
R989 vss.t85 vss.n103 5.2005
R990 vss.n1639 vss.n1638 5.2005
R991 vss.n1638 vss.n1637 5.2005
R992 vss.n168 vss.n167 5.2005
R993 vss.n168 vss.n97 5.2005
R994 vss.n115 vss.n110 5.2005
R995 vss.n1637 vss.n110 5.2005
R996 vss.n175 vss.n98 5.2005
R997 vss.t85 vss.n98 5.2005
R998 vss.n1644 vss.n99 5.2005
R999 vss.n1644 vss.n1643 5.2005
R1000 vss.n1647 vss.n1646 5.2005
R1001 vss.n1646 vss.n92 5.2005
R1002 vss.n96 vss.n94 5.2005
R1003 vss.n96 vss.t18 5.2005
R1004 vss.n1113 vss.n82 5.2005
R1005 vss.n1659 vss.n82 5.2005
R1006 vss.n1336 vss.n453 5.2005
R1007 vss.n1332 vss.n453 5.2005
R1008 vss.n1323 vss.n462 5.2005
R1009 vss.n1200 vss.n462 5.2005
R1010 vss.n1322 vss.n1321 5.2005
R1011 vss.n1321 vss.n457 5.2005
R1012 vss.n1328 vss.n452 5.2005
R1013 vss.n1331 vss.n452 5.2005
R1014 vss.n1329 vss.n1328 5.2005
R1015 vss.n1330 vss.n1329 5.2005
R1016 vss.n1351 vss.n1350 5.2005
R1017 vss.n1350 vss.n446 5.2005
R1018 vss.n1355 vss.n1354 5.2005
R1019 vss.n1356 vss.n1355 5.2005
R1020 vss.n1358 vss.n444 5.2005
R1021 vss.n1358 vss.n1357 5.2005
R1022 vss.n1335 vss.n1334 5.2005
R1023 vss.n1334 vss.n1333 5.2005
R1024 vss.n1390 vss.n438 5.2005
R1025 vss.n442 vss.n438 5.2005
R1026 vss.n1385 vss.n1384 5.2005
R1027 vss.n441 vss.n440 5.2005
R1028 vss.n1389 vss.n1388 5.2005
R1029 vss.n1388 vss.n1387 5.2005
R1030 vss.n1376 vss.n1363 5.2005
R1031 vss.n1366 vss.n1365 5.2005
R1032 vss.n1369 vss.n433 5.2005
R1033 vss.n433 vss.n401 5.2005
R1034 vss.n1375 vss.n1374 5.2005
R1035 vss.n1368 vss.n1367 5.2005
R1036 vss.n1371 vss.n1370 5.2005
R1037 vss.n1372 vss.n1371 5.2005
R1038 vss.n1115 vss.n1114 5.2005
R1039 vss.n1112 vss.n1110 5.2005
R1040 vss.n1197 vss.n1196 5.2005
R1041 vss.n1195 vss.n88 5.2005
R1042 vss.n1089 vss.n1088 5.2005
R1043 vss.n1093 vss.n1092 5.2005
R1044 vss.n1094 vss.n1093 5.2005
R1045 vss.n1090 vss.n1077 5.2005
R1046 vss.n1095 vss.n1077 5.2005
R1047 vss.n1107 vss.n1106 5.2005
R1048 vss.n1106 vss.n1105 5.2005
R1049 vss.n1103 vss.n1102 5.2005
R1050 vss.n1104 vss.n1103 5.2005
R1051 vss.n1100 vss.n1099 5.2005
R1052 vss.n1099 vss.n1074 5.2005
R1053 vss.n1097 vss.n1078 5.2005
R1054 vss.n1097 vss.n1096 5.2005
R1055 vss.n1086 vss.n1085 5.2005
R1056 vss.n330 vss.n325 5.2005
R1057 vss.n1501 vss.n1500 5.2005
R1058 vss.n1504 vss.n1503 5.2005
R1059 vss.n1507 vss.n1506 5.2005
R1060 vss.n1497 vss.n1491 5.2005
R1061 vss.n1510 vss.n330 5.2005
R1062 vss.n454 vss.n403 5.2005
R1063 vss.n407 vss.n403 5.2005
R1064 vss.n1442 vss.n404 5.2005
R1065 vss.n1442 vss.t0 5.2005
R1066 vss.n1443 vss.n352 5.2005
R1067 vss.t1 vss.n1443 5.2005
R1068 vss.n1489 vss.n350 5.2005
R1069 vss.n1460 vss.n350 5.2005
R1070 vss.n1520 vss.n1519 5.2005
R1071 vss.t9 vss.n1520 5.2005
R1072 vss.n1518 vss.n351 5.2005
R1073 vss.n351 vss.n335 5.2005
R1074 vss.n1486 vss.n355 5.2005
R1075 vss.n385 vss.n355 5.2005
R1076 vss.n1338 vss.n1337 5.2005
R1077 vss.n1340 vss.n451 5.2005
R1078 vss.n1344 vss.n1343 5.2005
R1079 vss.n1343 vss.n417 5.2005
R1080 vss.n1347 vss.n1346 5.2005
R1081 vss.n1349 vss.n448 5.2005
R1082 vss.n1352 vss.n447 5.2005
R1083 vss.n447 vss.n417 5.2005
R1084 vss.n1353 vss.n445 5.2005
R1085 vss.n445 vss.n417 5.2005
R1086 vss.n1360 vss.n1359 5.2005
R1087 vss.n1359 vss.n417 5.2005
R1088 vss.n1526 vss.n346 5.2005
R1089 vss.n346 vss.n335 5.2005
R1090 vss.n1524 vss.n345 5.2005
R1091 vss.t9 vss.n345 5.2005
R1092 vss.n348 vss.n347 5.2005
R1093 vss.n1460 vss.n348 5.2005
R1094 vss.n1447 vss.n395 5.2005
R1095 vss.t1 vss.n395 5.2005
R1096 vss.n397 vss.n396 5.2005
R1097 vss.t0 vss.n397 5.2005
R1098 vss.n1438 vss.n408 5.2005
R1099 vss.n408 vss.n407 5.2005
R1100 vss.n1615 vss.n208 5.2005
R1101 vss.n1615 vss.n1614 5.2005
R1102 vss.n1543 vss.n327 5.2005
R1103 vss.n1543 vss.n1542 5.2005
R1104 vss.n1525 vss.n326 5.2005
R1105 vss.n336 vss.n326 5.2005
R1106 vss.n1528 vss.n1527 5.2005
R1107 vss.n1529 vss.n1528 5.2005
R1108 vss.n1523 vss.n1522 5.2005
R1109 vss.n1522 vss.n1521 5.2005
R1110 vss.n388 vss.n387 5.2005
R1111 vss.n1461 vss.n388 5.2005
R1112 vss.n1474 vss.n1473 5.2005
R1113 vss.n1473 vss.n1472 5.2005
R1114 vss.n1477 vss.n1476 5.2005
R1115 vss.n1478 vss.n1477 5.2005
R1116 vss.n371 vss.n369 5.2005
R1117 vss.n369 vss.n357 5.2005
R1118 vss.n1449 vss.n1448 5.2005
R1119 vss.n1450 vss.n1449 5.2005
R1120 vss.n1446 vss.n1445 5.2005
R1121 vss.n1445 vss.n1444 5.2005
R1122 vss.n1440 vss.n1439 5.2005
R1123 vss.n1441 vss.n1440 5.2005
R1124 vss.n1437 vss.n1436 5.2005
R1125 vss.n1436 vss.n1435 5.2005
R1126 vss.n1361 vss.n409 5.2005
R1127 vss.n1420 vss.n409 5.2005
R1128 vss.n1382 vss.n1381 5.2005
R1129 vss.n1381 vss.n1380 5.2005
R1130 vss.n215 vss.n210 5.2005
R1131 vss.n1614 vss.n210 5.2005
R1132 vss.n341 vss.n329 5.2005
R1133 vss.n1542 vss.n329 5.2005
R1134 vss.n1532 vss.n1531 5.2005
R1135 vss.n1531 vss.n336 5.2005
R1136 vss.n1530 vss.n339 5.2005
R1137 vss.n1530 vss.n1529 5.2005
R1138 vss.n1465 vss.n343 5.2005
R1139 vss.n1521 vss.n343 5.2005
R1140 vss.n1468 vss.n1467 5.2005
R1141 vss.n1467 vss.n1461 5.2005
R1142 vss.n1463 vss.n367 5.2005
R1143 vss.n1472 vss.n367 5.2005
R1144 vss.n1480 vss.n1479 5.2005
R1145 vss.n1479 vss.n1478 5.2005
R1146 vss.n366 vss.n364 5.2005
R1147 vss.n366 vss.n357 5.2005
R1148 vss.n1426 vss.n394 5.2005
R1149 vss.n1450 vss.n394 5.2005
R1150 vss.n1428 vss.n399 5.2005
R1151 vss.n1444 vss.n399 5.2005
R1152 vss.n413 vss.n406 5.2005
R1153 vss.n1441 vss.n406 5.2005
R1154 vss.n1434 vss.n1433 5.2005
R1155 vss.n1435 vss.n1434 5.2005
R1156 vss.n415 vss.n411 5.2005
R1157 vss.n1420 vss.n411 5.2005
R1158 vss.n1379 vss.n1378 5.2005
R1159 vss.n1380 vss.n1379 5.2005
R1160 vss.n1612 vss.n1611 5.2005
R1161 vss.n1613 vss.n1612 5.2005
R1162 vss.n340 vss.n213 5.2005
R1163 vss.n213 vss.n209 5.2005
R1164 vss.n342 vss.n338 5.2005
R1165 vss.n338 vss.n328 5.2005
R1166 vss.n1534 vss.n1533 5.2005
R1167 vss.n1535 vss.n1534 5.2005
R1168 vss.n1464 vss.n337 5.2005
R1169 vss.n344 vss.n337 5.2005
R1170 vss.n1466 vss.n1462 5.2005
R1171 vss.n1462 vss.n349 5.2005
R1172 vss.n1470 vss.n1469 5.2005
R1173 vss.n1471 vss.n1470 5.2005
R1174 vss.n365 vss.n363 5.2005
R1175 vss.n368 vss.n363 5.2005
R1176 vss.n1482 vss.n1481 5.2005
R1177 vss.n1483 vss.n1482 5.2005
R1178 vss.n1425 vss.n362 5.2005
R1179 vss.n1451 vss.n362 5.2005
R1180 vss.n1427 vss.n1424 5.2005
R1181 vss.n1424 vss.n393 5.2005
R1182 vss.n1430 vss.n1429 5.2005
R1183 vss.n1430 vss.n398 5.2005
R1184 vss.n1432 vss.n1431 5.2005
R1185 vss.n1431 vss.n405 5.2005
R1186 vss.n1423 vss.n412 5.2005
R1187 vss.n1423 vss.n410 5.2005
R1188 vss.n1422 vss.n416 5.2005
R1189 vss.n1422 vss.n1421 5.2005
R1190 vss.n1377 vss.n414 5.2005
R1191 vss.n1362 vss.n414 5.2005
R1192 vss.n1594 vss.n225 5.2005
R1193 vss.n1594 vss.n1593 5.2005
R1194 vss.n332 vss.n211 5.2005
R1195 vss.n1613 vss.n211 5.2005
R1196 vss.n1539 vss.n1538 5.2005
R1197 vss.n1538 vss.n209 5.2005
R1198 vss.n1537 vss.n331 5.2005
R1199 vss.n1537 vss.n328 5.2005
R1200 vss.n1536 vss.n334 5.2005
R1201 vss.n1536 vss.n1535 5.2005
R1202 vss.n1456 vss.n333 5.2005
R1203 vss.n344 vss.n333 5.2005
R1204 vss.n1457 vss.n390 5.2005
R1205 vss.n390 vss.n349 5.2005
R1206 vss.n1459 vss.n1458 5.2005
R1207 vss.n1471 vss.n1459 5.2005
R1208 vss.n1455 vss.n389 5.2005
R1209 vss.n389 vss.n368 5.2005
R1210 vss.n1454 vss.n361 5.2005
R1211 vss.n1483 vss.n361 5.2005
R1212 vss.n1453 vss.n1452 5.2005
R1213 vss.n1452 vss.n1451 5.2005
R1214 vss.n392 vss.n391 5.2005
R1215 vss.n393 vss.n392 5.2005
R1216 vss.n1414 vss.n1413 5.2005
R1217 vss.n1414 vss.n398 5.2005
R1218 vss.n1416 vss.n1415 5.2005
R1219 vss.n1415 vss.n405 5.2005
R1220 vss.n1417 vss.n419 5.2005
R1221 vss.n419 vss.n410 5.2005
R1222 vss.n1419 vss.n1418 5.2005
R1223 vss.n1421 vss.n1419 5.2005
R1224 vss.n1409 vss.n418 5.2005
R1225 vss.n1362 vss.n418 5.2005
R1226 vss.n1408 vss.n1407 5.2005
R1227 vss.n422 vss.n421 5.2005
R1228 vss.n1404 vss.n1403 5.2005
R1229 vss.n1405 vss.n1404 5.2005
R1230 vss.n741 vss.n740 5.2005
R1231 vss.n747 vss.n746 5.2005
R1232 vss.n748 vss.n742 5.2005
R1233 vss.n744 vss.n742 5.2005
R1234 vss.n776 vss.n775 5.2005
R1235 vss.n775 vss.n737 5.2005
R1236 vss.n781 vss.n780 5.2005
R1237 vss.n773 vss.n739 5.2005
R1238 vss.n750 vss.n736 5.2005
R1239 vss.n792 vss.n736 5.2005
R1240 vss.n751 vss.n743 5.2005
R1241 vss.n743 vss.t5 5.2005
R1242 vss.n753 vss.n752 5.2005
R1243 vss.n754 vss.n753 5.2005
R1244 vss.n756 vss.n755 5.2005
R1245 vss.n755 vss.n754 5.2005
R1246 vss.n757 vss.n738 5.2005
R1247 vss.n738 vss.t5 5.2005
R1248 vss.n791 vss.n790 5.2005
R1249 vss.n792 vss.n791 5.2005
R1250 vss.n765 vss.n764 5.2005
R1251 vss.n766 vss.n763 5.2005
R1252 vss.n768 vss.n767 5.2005
R1253 vss.n769 vss.n768 5.2005
R1254 vss.n760 vss.n759 5.2005
R1255 vss.n770 vss.n760 5.2005
R1256 vss.n788 vss.n787 5.2005
R1257 vss.n787 vss.n786 5.2005
R1258 vss.n774 vss.n679 5.2005
R1259 vss.n680 vss.n679 5.2005
R1260 vss.n778 vss.n777 5.2005
R1261 vss.n777 vss.n771 5.2005
R1262 vss.n783 vss.n782 5.2005
R1263 vss.n784 vss.n783 5.2005
R1264 vss.n761 vss.n758 5.2005
R1265 vss.n785 vss.n761 5.2005
R1266 vss.n803 vss.n678 5.2005
R1267 vss.n803 vss.n802 5.2005
R1268 vss.n834 vss.n629 5.2005
R1269 vss.n835 vss.n834 5.2005
R1270 vss.n833 vss.n832 5.2005
R1271 vss.n833 vss.t54 5.2005
R1272 vss.n831 vss.n662 5.2005
R1273 vss.n673 vss.n662 5.2005
R1274 vss.n829 vss.n828 5.2005
R1275 vss.n828 vss.n827 5.2005
R1276 vss.n665 vss.n664 5.2005
R1277 vss.t58 vss.n665 5.2005
R1278 vss.n825 vss.n672 5.2005
R1279 vss.n825 vss.n824 5.2005
R1280 vss.n648 vss.n637 5.2005
R1281 vss.n645 vss.n644 5.2005
R1282 vss.n645 vss.n545 5.2005
R1283 vss.n642 vss.n641 5.2005
R1284 vss.n639 vss.n638 5.2005
R1285 vss.n651 vss.n650 5.2005
R1286 vss.n653 vss.n635 5.2005
R1287 vss.n635 vss.n545 5.2005
R1288 vss.n841 vss.n636 5.2005
R1289 vss.n636 vss.n545 5.2005
R1290 vss.n839 vss.n838 5.2005
R1291 vss.n838 vss.n545 5.2005
R1292 vss.n836 vss.n661 5.2005
R1293 vss.n836 vss.n835 5.2005
R1294 vss.n807 vss.n660 5.2005
R1295 vss.t54 vss.n660 5.2005
R1296 vss.n810 vss.n809 5.2005
R1297 vss.n809 vss.n673 5.2005
R1298 vss.n806 vss.n667 5.2005
R1299 vss.n827 vss.n667 5.2005
R1300 vss.n805 vss.n804 5.2005
R1301 vss.n804 vss.t58 5.2005
R1302 vss.n909 vss.n908 5.2005
R1303 vss.n910 vss.n909 5.2005
R1304 vss.n907 vss.n550 5.2005
R1305 vss.n550 vss.n548 5.2005
R1306 vss.n919 vss.n918 5.2005
R1307 vss.n920 vss.n919 5.2005
R1308 vss.n914 vss.n549 5.2005
R1309 vss.n920 vss.n549 5.2005
R1310 vss.n913 vss.n912 5.2005
R1311 vss.n912 vss.n548 5.2005
R1312 vss.n911 vss.n553 5.2005
R1313 vss.n911 vss.n910 5.2005
R1314 vss.n916 vss.n915 5.2005
R1315 vss.n917 vss.n551 5.2005
R1316 vss.n892 vss.n891 5.2005
R1317 vss.n891 vss.n890 5.2005
R1318 vss.n617 vss.n616 5.2005
R1319 vss.t3 vss.n617 5.2005
R1320 vss.n851 vss.n850 5.2005
R1321 vss.n852 vss.n851 5.2005
R1322 vss.n849 vss.n628 5.2005
R1323 vss.n844 vss.n628 5.2005
R1324 vss.n847 vss.n846 5.2005
R1325 vss.n876 vss.n557 5.2005
R1326 vss.n879 vss.n878 5.2005
R1327 vss.n874 vss.n622 5.2005
R1328 vss.n622 vss.n559 5.2005
R1329 vss.n627 vss.n623 5.2005
R1330 vss.n852 vss.n627 5.2005
R1331 vss.n855 vss.n621 5.2005
R1332 vss.n621 vss.t3 5.2005
R1333 vss.n889 vss.n888 5.2005
R1334 vss.n890 vss.n889 5.2005
R1335 vss.n853 vss.n623 5.2005
R1336 vss.n853 vss.n852 5.2005
R1337 vss.n855 vss.n854 5.2005
R1338 vss.n854 vss.t3 5.2005
R1339 vss.n888 vss.n619 5.2005
R1340 vss.n890 vss.n619 5.2005
R1341 vss.n632 vss.n630 5.2005
R1342 vss.n868 vss.n867 5.2005
R1343 vss.n865 vss.n864 5.2005
R1344 vss.n860 vss.n618 5.2005
R1345 vss.n618 vss.n559 5.2005
R1346 vss.n652 vss.n633 5.2005
R1347 vss.n844 vss.n633 5.2005
R1348 vss.n843 vss.n842 5.2005
R1349 vss.n844 vss.n843 5.2005
R1350 vss.n840 vss.n634 5.2005
R1351 vss.n844 vss.n634 5.2005
R1352 vss.n654 vss.n620 5.2005
R1353 vss.n890 vss.n620 5.2005
R1354 vss.n656 vss.n655 5.2005
R1355 vss.n655 vss.t3 5.2005
R1356 vss.n657 vss.n626 5.2005
R1357 vss.n852 vss.n626 5.2005
R1358 vss.n613 vss.n612 5.2005
R1359 vss.n612 vss.n611 5.2005
R1360 vss.n614 vss.n569 5.2005
R1361 vss.n569 vss.n566 5.2005
R1362 vss.n900 vss.n899 5.2005
R1363 vss.n898 vss.n568 5.2005
R1364 vss.n897 vss.n567 5.2005
R1365 vss.n902 vss.n567 5.2005
R1366 vss.n896 vss.n895 5.2005
R1367 vss.n857 vss.n615 5.2005
R1368 vss.n859 vss.n858 5.2005
R1369 vss.n863 vss.n862 5.2005
R1370 vss.n861 vss.n856 5.2005
R1371 vss.n870 vss.n869 5.2005
R1372 vss.n872 vss.n871 5.2005
R1373 vss.n884 vss.n873 5.2005
R1374 vss.n886 vss.n885 5.2005
R1375 vss.n883 vss.n882 5.2005
R1376 vss.n881 vss.n880 5.2005
R1377 vss.n875 vss.n558 5.2005
R1378 vss.n905 vss.n904 5.2005
R1379 vss.n906 vss.n556 5.2005
R1380 vss.n575 vss.n554 5.2005
R1381 vss.n577 vss.n576 5.2005
R1382 vss.n579 vss.n578 5.2005
R1383 vss.n580 vss.n574 5.2005
R1384 vss.n582 vss.n581 5.2005
R1385 vss.n591 vss.n541 5.2005
R1386 vss.n593 vss.n592 5.2005
R1387 vss.n595 vss.n594 5.2005
R1388 vss.n597 vss.n596 5.2005
R1389 vss.n599 vss.n598 5.2005
R1390 vss.n601 vss.n600 5.2005
R1391 vss.n603 vss.n602 5.2005
R1392 vss.n605 vss.n604 5.2005
R1393 vss.n606 vss.n589 5.2005
R1394 vss.n608 vss.n607 5.2005
R1395 vss.n590 vss.n588 5.2005
R1396 vss.n571 vss.n570 5.2005
R1397 vss.n610 vss.n571 5.2005
R1398 vss.n711 vss.n710 5.2005
R1399 vss.n710 vss.n547 5.2005
R1400 vss.n706 vss.n705 5.2005
R1401 vss.n708 vss.n701 5.2005
R1402 vss.n709 vss.n700 5.2005
R1403 vss.n709 vss.n625 5.2005
R1404 vss.n703 vss.n702 5.2005
R1405 vss.n702 vss.n547 5.2005
R1406 vss.n1285 vss.n1284 5.2005
R1407 vss.n1286 vss.n1285 5.2005
R1408 vss.n1275 vss.n511 5.2005
R1409 vss.n1211 vss.n511 5.2005
R1410 vss.n1274 vss.n1273 5.2005
R1411 vss.n1271 vss.n513 5.2005
R1412 vss.n1270 vss.n1269 5.2005
R1413 vss.n1270 vss.n6 5.2005
R1414 vss.n1268 vss.n514 5.2005
R1415 vss.n1267 vss.n1266 5.2005
R1416 vss.n1264 vss.n515 5.2005
R1417 vss.n1262 vss.n1261 5.2005
R1418 vss.n1260 vss.n516 5.2005
R1419 vss.n1259 vss.n1258 5.2005
R1420 vss.n1256 vss.n517 5.2005
R1421 vss.n1254 vss.n1253 5.2005
R1422 vss.n1252 vss.n518 5.2005
R1423 vss.n1251 vss.n1250 5.2005
R1424 vss.n1248 vss.n519 5.2005
R1425 vss.n1246 vss.n1245 5.2005
R1426 vss.n1244 vss.n520 5.2005
R1427 vss.n1243 vss.n1242 5.2005
R1428 vss.n1240 vss.n521 5.2005
R1429 vss.n1238 vss.n1237 5.2005
R1430 vss.n1236 vss.n522 5.2005
R1431 vss.n522 vss.n6 5.2005
R1432 vss.n1287 vss.n508 5.2005
R1433 vss.n1287 vss.n1286 5.2005
R1434 vss.n523 vss.n507 5.2005
R1435 vss.n1211 vss.n507 5.2005
R1436 vss.n1309 vss.n1308 5.2005
R1437 vss.n471 vss.n469 5.2005
R1438 vss.n1305 vss.n1304 5.2005
R1439 vss.n1306 vss.n1305 5.2005
R1440 vss.n1320 vss.n461 5.2005
R1441 vss.n461 vss.n426 5.2005
R1442 vss.n1325 vss.n1324 5.2005
R1443 vss.t37 vss.n1325 5.2005
R1444 vss.n1327 vss.n1326 5.2005
R1445 vss.n1326 vss.t37 5.2005
R1446 vss.n460 vss.n459 5.2005
R1447 vss.n460 vss.n426 5.2005
R1448 vss.n1327 vss.n458 5.2005
R1449 vss.t37 vss.n458 5.2005
R1450 vss.n496 vss.n459 5.2005
R1451 vss.n496 vss.n426 5.2005
R1452 vss.n498 vss.n497 5.2005
R1453 vss.n501 vss.n500 5.2005
R1454 vss.n481 vss.n474 5.2005
R1455 vss.n1306 vss.n474 5.2005
R1456 vss.n439 vss.n437 5.2005
R1457 vss.t37 vss.n437 5.2005
R1458 vss.n1299 vss.n1298 5.2005
R1459 vss.n1298 vss.n426 5.2005
R1460 vss.n1294 vss.n1293 5.2005
R1461 vss.n503 vss.n502 5.2005
R1462 vss.n499 vss.n482 5.2005
R1463 vss.n495 vss.n494 5.2005
R1464 vss.n492 vss.n483 5.2005
R1465 vss.n490 vss.n489 5.2005
R1466 vss.n487 vss.n486 5.2005
R1467 vss.n484 vss.n470 5.2005
R1468 vss.n1311 vss.n1310 5.2005
R1469 vss.n1313 vss.n467 5.2005
R1470 vss.n1314 vss.n464 5.2005
R1471 vss.n1317 vss.n1316 5.2005
R1472 vss.n465 vss.n463 5.2005
R1473 vss.n1279 vss.n1277 5.2005
R1474 vss.n1280 vss.n1276 5.2005
R1475 vss.n1283 vss.n1282 5.2005
R1476 vss.n1289 vss.n505 5.2005
R1477 vss.n506 vss.n505 5.2005
R1478 vss.n506 vss.n466 5.2005
R1479 vss.n1292 vss.n466 5.2005
R1480 vss.n1392 vss.n1391 5.2005
R1481 vss.n1393 vss.n1392 5.2005
R1482 vss.n1297 vss.n1296 5.2005
R1483 vss.n1297 vss.n427 5.2005
R1484 vss.n1300 vss.n479 5.2005
R1485 vss.n479 vss.n478 5.2005
R1486 vss.n1302 vss.n1301 5.2005
R1487 vss.n1303 vss.n1302 5.2005
R1488 vss.n1216 vss.n480 5.2005
R1489 vss.n1216 vss.n63 5.2005
R1490 vss.n1219 vss.n1218 5.2005
R1491 vss.n1220 vss.n1219 5.2005
R1492 vss.n1217 vss.n1214 5.2005
R1493 vss.n1214 vss.n510 5.2005
R1494 vss.n1213 vss.n1210 5.2005
R1495 vss.n1213 vss.n1212 5.2005
R1496 vss.n1234 vss.n1233 5.2005
R1497 vss.n527 vss.n524 5.2005
R1498 vss.n1230 vss.n1229 5.2005
R1499 vss.n1231 vss.n1230 5.2005
R1500 vss.n1394 vss.n434 5.2005
R1501 vss.n1394 vss.n1393 5.2005
R1502 vss.n1396 vss.n1395 5.2005
R1503 vss.n1395 vss.n427 5.2005
R1504 vss.n432 vss.n430 5.2005
R1505 vss.n478 vss.n432 5.2005
R1506 vss.n1049 vss.n475 5.2005
R1507 vss.n1303 vss.n475 5.2005
R1508 vss.n1051 vss.n537 5.2005
R1509 vss.n537 vss.n63 5.2005
R1510 vss.n1221 vss.n538 5.2005
R1511 vss.n1221 vss.n1220 5.2005
R1512 vss.n1223 vss.n1222 5.2005
R1513 vss.n1222 vss.n510 5.2005
R1514 vss.n536 vss.n532 5.2005
R1515 vss.n1212 vss.n536 5.2005
R1516 vss.n431 vss.n429 5.2005
R1517 vss.n435 vss.n429 5.2005
R1518 vss.n1398 vss.n1397 5.2005
R1519 vss.n1399 vss.n1398 5.2005
R1520 vss.n1048 vss.n428 5.2005
R1521 vss.n477 vss.n428 5.2005
R1522 vss.n1050 vss.n1047 5.2005
R1523 vss.n1047 vss.n472 5.2005
R1524 vss.n1053 vss.n1052 5.2005
R1525 vss.n1054 vss.n1053 5.2005
R1526 vss.n535 vss.n534 5.2005
R1527 vss.n1063 vss.n534 5.2005
R1528 vss.n1225 vss.n1224 5.2005
R1529 vss.n1225 vss.n509 5.2005
R1530 vss.n1227 vss.n1226 5.2005
R1531 vss.n1226 vss.n529 5.2005
R1532 vss.n1041 vss.n531 5.2005
R1533 vss.n1043 vss.n1039 5.2005
R1534 vss.n1402 vss.n423 5.2005
R1535 vss.n435 vss.n423 5.2005
R1536 vss.n1401 vss.n1400 5.2005
R1537 vss.n1400 vss.n1399 5.2005
R1538 vss.n425 vss.n424 5.2005
R1539 vss.n477 vss.n425 5.2005
R1540 vss.n1058 vss.n1057 5.2005
R1541 vss.n1057 vss.n472 5.2005
R1542 vss.n1060 vss.n540 5.2005
R1543 vss.n1054 vss.n540 5.2005
R1544 vss.n1062 vss.n1061 5.2005
R1545 vss.n1063 vss.n1062 5.2005
R1546 vss.n1046 vss.n539 5.2005
R1547 vss.n539 vss.n509 5.2005
R1548 vss.n1045 vss.n1044 5.2005
R1549 vss.n1044 vss.n529 5.2005
R1550 vss.n1204 vss.n1203 5.2005
R1551 vss.n1203 vss.n1202 5.2005
R1552 vss.n1068 vss.n1066 5.2005
R1553 vss.n1066 vss.n66 5.2005
R1554 vss.n1209 vss.n1208 5.2005
R1555 vss.t76 vss.n1209 5.2005
R1556 vss.n1067 vss.n1065 5.2005
R1557 vss.n1180 vss.n1065 5.2005
R1558 vss.n1124 vss.n1123 5.2005
R1559 vss.n1194 vss.n1111 5.2005
R1560 vss.n1202 vss.n1111 5.2005
R1561 vss.n1192 vss.n1191 5.2005
R1562 vss.n1191 vss.n66 5.2005
R1563 vss.n1183 vss.n1064 5.2005
R1564 vss.t76 vss.n1064 5.2005
R1565 vss.n1182 vss.n1181 5.2005
R1566 vss.n1181 vss.n1180 5.2005
R1567 vss.n1189 vss.n1118 5.2005
R1568 vss.n1187 vss.n1186 5.2005
R1569 vss.n1185 vss.n1184 5.2005
R1570 vss.n1184 vss.n75 5.2005
R1571 vss.n1665 vss.n1664 5.2005
R1572 vss.n1666 vss.n1665 5.2005
R1573 vss.n62 vss.n60 5.2005
R1574 vss.t27 vss.n62 5.2005
R1575 vss.n1674 vss.n1673 5.2005
R1576 vss.n1673 vss.n1672 5.2005
R1577 vss.n1133 vss.n61 5.2005
R1578 vss.n1177 vss.n1176 5.2005
R1579 vss.n1131 vss.n1129 5.2005
R1580 vss.n1179 vss.n1129 5.2005
R1581 vss.n1668 vss.n71 5.2005
R1582 vss.n1666 vss.n71 5.2005
R1583 vss.n1669 vss.n70 5.2005
R1584 vss.t27 vss.n70 5.2005
R1585 vss.n1670 vss.n64 5.2005
R1586 vss.n1672 vss.n64 5.2005
R1587 vss.n1668 vss.n1667 5.2005
R1588 vss.n1667 vss.n1666 5.2005
R1589 vss.n1669 vss.n68 5.2005
R1590 vss.t27 vss.n68 5.2005
R1591 vss.n1671 vss.n1670 5.2005
R1592 vss.n1672 vss.n1671 5.2005
R1593 vss.n1163 vss.n67 5.2005
R1594 vss.n1141 vss.n1140 5.2005
R1595 vss.n1145 vss.n1128 5.2005
R1596 vss.n1179 vss.n1128 5.2005
R1597 vss.n1098 vss.n1076 5.2005
R1598 vss.n1098 vss.n436 5.2005
R1599 vss.n1101 vss.n1075 5.2005
R1600 vss.n1075 vss.n436 5.2005
R1601 vss.n1072 vss.n1071 5.2005
R1602 vss.n1072 vss.n436 5.2005
R1603 vss.n1663 vss.n76 5.2005
R1604 vss.n436 vss.n76 5.2005
R1605 vss.n1084 vss.n1081 5.2005
R1606 vss.n1082 vss.n77 5.2005
R1607 vss.n1666 vss.n74 5.2005
R1608 vss.n1153 vss.t27 5.2005
R1609 vss.n1155 vss.n65 5.2005
R1610 vss.n1672 vss.n65 5.2005
R1611 vss.n54 vss.n7 5.2005
R1612 vss.n53 vss.n52 5.2005
R1613 vss.n50 vss.n9 5.2005
R1614 vss.n50 vss.n5 5.2005
R1615 vss.n49 vss.n48 5.2005
R1616 vss.n47 vss.n46 5.2005
R1617 vss.n45 vss.n11 5.2005
R1618 vss.n43 vss.n42 5.2005
R1619 vss.n41 vss.n12 5.2005
R1620 vss.n40 vss.n39 5.2005
R1621 vss.n37 vss.n13 5.2005
R1622 vss.n35 vss.n34 5.2005
R1623 vss.n33 vss.n14 5.2005
R1624 vss.n32 vss.n31 5.2005
R1625 vss.n29 vss.n15 5.2005
R1626 vss.n27 vss.n26 5.2005
R1627 vss.n25 vss.n16 5.2005
R1628 vss.n24 vss.n23 5.2005
R1629 vss.n21 vss.n17 5.2005
R1630 vss.n19 vss.n18 5.2005
R1631 vss.n3 vss.n1 5.2005
R1632 vss.n5 vss.n3 5.2005
R1633 vss.n1148 vss.n1070 5.2005
R1634 vss.n1150 vss.n1146 5.2005
R1635 vss.n1152 vss.n1151 5.2005
R1636 vss.n1156 vss.n1144 5.2005
R1637 vss.n1158 vss.n1157 5.2005
R1638 vss.n1160 vss.n1143 5.2005
R1639 vss.n1162 vss.n1161 5.2005
R1640 vss.n1164 vss.n1139 5.2005
R1641 vss.n1166 vss.n1165 5.2005
R1642 vss.n1169 vss.n1168 5.2005
R1643 vss.n1171 vss.n1170 5.2005
R1644 vss.n1173 vss.n1138 5.2005
R1645 vss.n1175 vss.n1174 5.2005
R1646 vss.n1136 vss.n1130 5.2005
R1647 vss.n1135 vss.n1134 5.2005
R1648 vss.n59 vss.n58 5.2005
R1649 vss.n1678 vss.n1677 5.2005
R1650 vss.n1680 vss.n57 5.2005
R1651 vss.n1681 vss.n55 5.2005
R1652 vss.n1684 vss.n1683 5.2005
R1653 vss.n4 vss.n2 5.2005
R1654 vss.n528 vss.n4 5.2005
R1655 vss.n1690 vss.n1689 5.2005
R1656 vss.n1689 vss.n1688 5.2005
R1657 vss.n1687 vss.n1686 5.2005
R1658 vss.n1688 vss.n1687 5.2005
R1659 vss.n1685 vss.n8 5.2005
R1660 vss.n528 vss.n8 5.2005
R1661 vss.n712 vss.n699 5.2005
R1662 vss.n699 vss.n546 5.2005
R1663 vss.n714 vss.n713 5.2005
R1664 vss.n715 vss.n714 5.2005
R1665 vss.n693 vss.n691 5.2005
R1666 vss.n695 vss.n693 5.2005
R1667 vss.n724 vss.n723 5.2005
R1668 vss.n694 vss.n692 5.2005
R1669 vss.n720 vss.n719 5.2005
R1670 vss.n721 vss.n720 5.2005
R1671 vss.n698 vss.n697 5.2005
R1672 vss.n698 vss.n546 5.2005
R1673 vss.n717 vss.n716 5.2005
R1674 vss.n716 vss.n715 5.2005
R1675 vss.n718 vss.n696 5.2005
R1676 vss.n696 vss.n695 5.2005
R1677 vss.n780 vss.n772 5.15839
R1678 vss.n484 vss.n468 4.98535
R1679 vss.n1499 vss.n1498 4.93742
R1680 vss.n1496 vss.n1490 4.93742
R1681 vss.n631 vss.n628 4.61478
R1682 vss.n79 vss.n76 4.61478
R1683 vss.n1321 vss.n456 4.61478
R1684 vss.n1460 vss.n349 4.59479
R1685 vss.t9 vss.n344 4.59479
R1686 vss.n1535 vss.n335 4.59479
R1687 vss.n1591 vss.n224 4.46256
R1688 vss.t10 vss.n1590 4.46256
R1689 vss.n1231 vss.n528 4.46256
R1690 vss.n1615 vss.n206 4.27828
R1691 vss.n775 vss.n772 4.23734
R1692 vss.n824 vss.n666 4.17792
R1693 vss.n808 vss.n672 4.17792
R1694 vss.n167 vss.n102 4.04738
R1695 vss.n1645 vss.n97 4.04738
R1696 vss.n1486 vss.n354 4.04738
R1697 vss.n187 vss.n148 3.8757
R1698 vss.n838 vss.n837 3.62288
R1699 vss.n1106 vss.n1073 3.62288
R1700 vss.n1291 vss.n1290 3.61637
R1701 vss.n1561 vss.n232 3.51433
R1702 vss.n787 vss.n761 3.38837
R1703 vss.n1547 vss.n323 3.35907
R1704 vss.n1617 vss.n204 3.24563
R1705 vss.n233 vss.n229 3.24563
R1706 vss.n1180 vss.n1179 3.24563
R1707 vss.n1666 vss.n75 3.24563
R1708 vss.n1202 vss.n436 3.24563
R1709 vss.n1562 vss.n227 3.21767
R1710 vss.n1288 vss.n506 3.08259
R1711 vss.n385 vss.n370 3.00831
R1712 vss.n1359 vss.n443 2.69281
R1713 vss.n1281 vss.n1280 2.65224
R1714 vss.n1278 vss.n465 2.65224
R1715 vss.n1315 vss.n1314 2.65224
R1716 vss.n1312 vss.n1311 2.65224
R1717 vss.n486 vss.n485 2.65224
R1718 vss.n492 vss.n491 2.65224
R1719 vss.n493 vss.n482 2.65224
R1720 vss.n1293 vss.n504 2.65224
R1721 vss.n504 vss.n503 2.65224
R1722 vss.n494 vss.n493 2.65224
R1723 vss.n491 vss.n490 2.65224
R1724 vss.n485 vss.n484 2.65224
R1725 vss.n1313 vss.n1312 2.65224
R1726 vss.n1316 vss.n1315 2.65224
R1727 vss.n1279 vss.n1278 2.65224
R1728 vss.n1282 vss.n1281 2.65224
R1729 vss.n167 vss.n166 2.6005
R1730 vss.n165 vss.n164 2.6005
R1731 vss.n163 vss.n162 2.6005
R1732 vss.n160 vss.n159 2.6005
R1733 vss.n158 vss.n157 2.6005
R1734 vss.n152 vss.n151 2.6005
R1735 vss.n172 vss.n171 2.6005
R1736 vss.n173 vss.n97 2.6005
R1737 vss.n1487 vss.n1486 2.6005
R1738 vss.n356 vss.n353 2.6005
R1739 vss.n374 vss.n373 2.6005
R1740 vss.n376 vss.n375 2.6005
R1741 vss.n379 vss.n378 2.6005
R1742 vss.n381 vss.n380 2.6005
R1743 vss.n384 vss.n383 2.6005
R1744 vss.n386 vss.n385 2.6005
R1745 vss.n812 vss.n672 2.6005
R1746 vss.n814 vss.n813 2.6005
R1747 vss.n816 vss.n815 2.6005
R1748 vss.n818 vss.n817 2.6005
R1749 vss.n820 vss.n819 2.6005
R1750 vss.n822 vss.n821 2.6005
R1751 vss.n677 vss.n676 2.6005
R1752 vss.n824 vss.n663 2.6005
R1753 vss.n783 vss.n761 2.58746
R1754 vss.n777 vss.n679 2.58746
R1755 vss.n1659 vss.n1658 2.58397
R1756 vss.n783 vss.n772 2.51137
R1757 vss.n1097 vss.n1077 2.497
R1758 vss.n1334 vss.n453 2.497
R1759 vss.n1219 vss.n1216 2.48734
R1760 vss.n1085 vss.n1079 2.48287
R1761 vss.n1682 vss.n1681 2.46896
R1762 vss.n1679 vss.n1678 2.46896
R1763 vss.n1135 vss.n1132 2.46896
R1764 vss.n1174 vss.n1137 2.46896
R1765 vss.n1172 vss.n1171 2.46896
R1766 vss.n1167 vss.n1166 2.46896
R1767 vss.n1161 vss.n1142 2.46896
R1768 vss.n1159 vss.n1158 2.46896
R1769 vss.n1151 vss.n1147 2.46896
R1770 vss.n1149 vss.n1148 2.46896
R1771 vss.n51 vss.n7 2.46896
R1772 vss.n49 vss.n10 2.46896
R1773 vss.n45 vss.n44 2.46896
R1774 vss.n38 vss.n12 2.46896
R1775 vss.n37 vss.n36 2.46896
R1776 vss.n30 vss.n14 2.46896
R1777 vss.n29 vss.n28 2.46896
R1778 vss.n22 vss.n16 2.46896
R1779 vss.n21 vss.n20 2.46896
R1780 vss.n707 vss.n706 2.46896
R1781 vss.n723 vss.n722 2.46896
R1782 vss.n609 vss.n608 2.46896
R1783 vss.n604 vss.n587 2.46896
R1784 vss.n600 vss.n586 2.46896
R1785 vss.n596 vss.n585 2.46896
R1786 vss.n592 vss.n584 2.46896
R1787 vss.n583 vss.n582 2.46896
R1788 vss.n578 vss.n573 2.46896
R1789 vss.n572 vss.n554 2.46896
R1790 vss.n915 vss.n544 2.46896
R1791 vss.n901 vss.n900 2.46896
R1792 vss.n895 vss.n560 2.46896
R1793 vss.n858 vss.n561 2.46896
R1794 vss.n861 vss.n562 2.46896
R1795 vss.n871 vss.n563 2.46896
R1796 vss.n885 vss.n564 2.46896
R1797 vss.n881 vss.n565 2.46896
R1798 vss.n904 vss.n903 2.46896
R1799 vss.n992 vss.n972 2.46896
R1800 vss.n988 vss.n973 2.46896
R1801 vss.n978 vss.n963 2.46896
R1802 vss.n981 vss.n980 2.46896
R1803 vss.n956 vss.n936 2.46896
R1804 vss.n952 vss.n937 2.46896
R1805 vss.n942 vss.n927 2.46896
R1806 vss.n945 vss.n944 2.46896
R1807 vss.n942 vss.n941 2.46896
R1808 vss.n944 vss.n939 2.46896
R1809 vss.n955 vss.n937 2.46896
R1810 vss.n936 vss.n934 2.46896
R1811 vss.n978 vss.n977 2.46896
R1812 vss.n980 vss.n975 2.46896
R1813 vss.n991 vss.n973 2.46896
R1814 vss.n972 vss.n970 2.46896
R1815 vss.n877 vss.n876 2.46896
R1816 vss.n867 vss.n866 2.46896
R1817 vss.n780 vss.n779 2.46896
R1818 vss.n745 vss.n741 2.46896
R1819 vss.n1178 vss.n61 2.46896
R1820 vss.n1154 vss.n74 2.46896
R1821 vss.n1127 vss.n67 2.46896
R1822 vss.n126 vss.n121 2.46896
R1823 vss.n130 vss.n122 2.46896
R1824 vss.n124 vss.n123 2.46896
R1825 vss.n137 vss.n136 2.46896
R1826 vss.n302 vss.n301 2.46896
R1827 vss.n288 vss.n287 2.46896
R1828 vss.n278 vss.n265 2.46896
R1829 vss.n1116 vss.n1115 2.46896
R1830 vss.n1125 vss.n1124 2.46896
R1831 vss.n1189 vss.n1188 2.46896
R1832 vss.n1198 vss.n1197 2.46896
R1833 vss.n1653 vss.n83 2.46896
R1834 vss.n193 vss.n144 2.46896
R1835 vss.n1374 vss.n1373 2.46896
R1836 vss.n1364 vss.n1363 2.46896
R1837 vss.n1577 vss.n1576 2.46896
R1838 vss.n1509 vss.n1493 2.46896
R1839 vss.n1308 vss.n1307 2.46896
R1840 vss.n497 vss.n473 2.46896
R1841 vss.n1510 vss.n1490 2.46896
R1842 vss.n1497 vss.n1496 2.46896
R1843 vss.n1505 vss.n1504 2.46896
R1844 vss.n1498 vss.n325 2.46896
R1845 vss.n1273 vss.n1272 2.46896
R1846 vss.n1265 vss.n514 2.46896
R1847 vss.n1264 vss.n1263 2.46896
R1848 vss.n1257 vss.n516 2.46896
R1849 vss.n1256 vss.n1255 2.46896
R1850 vss.n1249 vss.n518 2.46896
R1851 vss.n1248 vss.n1247 2.46896
R1852 vss.n1241 vss.n520 2.46896
R1853 vss.n1240 vss.n1239 2.46896
R1854 vss.n1407 vss.n1406 2.46896
R1855 vss.n1567 vss.n1566 2.46896
R1856 vss.n1494 vss.n1493 2.46896
R1857 vss.n1578 vss.n1577 2.46896
R1858 vss.n1568 vss.n1567 2.46896
R1859 vss.n275 vss.n265 2.46896
R1860 vss.n302 vss.n260 2.46896
R1861 vss.n289 vss.n288 2.46896
R1862 vss.n85 vss.n83 2.46896
R1863 vss.n179 vss.n144 2.46896
R1864 vss.n137 vss.n135 2.46896
R1865 vss.n131 vss.n123 2.46896
R1866 vss.n127 vss.n122 2.46896
R1867 vss.n121 vss.n108 2.46896
R1868 vss.n1365 vss.n1364 2.46896
R1869 vss.n1373 vss.n1367 2.46896
R1870 vss.n1116 vss.n1110 2.46896
R1871 vss.n1198 vss.n88 2.46896
R1872 vss.n1500 vss.n1499 2.46896
R1873 vss.n1506 vss.n1505 2.46896
R1874 vss.n1406 vss.n422 2.46896
R1875 vss.n746 vss.n745 2.46896
R1876 vss.n779 vss.n739 2.46896
R1877 vss.n551 vss.n544 2.46896
R1878 vss.n878 vss.n877 2.46896
R1879 vss.n866 vss.n865 2.46896
R1880 vss.n901 vss.n568 2.46896
R1881 vss.n857 vss.n560 2.46896
R1882 vss.n862 vss.n561 2.46896
R1883 vss.n870 vss.n562 2.46896
R1884 vss.n884 vss.n563 2.46896
R1885 vss.n882 vss.n564 2.46896
R1886 vss.n565 vss.n558 2.46896
R1887 vss.n903 vss.n556 2.46896
R1888 vss.n577 vss.n572 2.46896
R1889 vss.n574 vss.n573 2.46896
R1890 vss.n591 vss.n583 2.46896
R1891 vss.n595 vss.n584 2.46896
R1892 vss.n599 vss.n585 2.46896
R1893 vss.n603 vss.n586 2.46896
R1894 vss.n589 vss.n587 2.46896
R1895 vss.n609 vss.n588 2.46896
R1896 vss.n708 vss.n707 2.46896
R1897 vss.n1272 vss.n1271 2.46896
R1898 vss.n1266 vss.n1265 2.46896
R1899 vss.n1263 vss.n1262 2.46896
R1900 vss.n1258 vss.n1257 2.46896
R1901 vss.n1255 vss.n1254 2.46896
R1902 vss.n1250 vss.n1249 2.46896
R1903 vss.n1247 vss.n1246 2.46896
R1904 vss.n1242 vss.n1241 2.46896
R1905 vss.n1239 vss.n1238 2.46896
R1906 vss.n1307 vss.n471 2.46896
R1907 vss.n500 vss.n473 2.46896
R1908 vss.n1126 vss.n1125 2.46896
R1909 vss.n1188 vss.n1187 2.46896
R1910 vss.n1178 vss.n1177 2.46896
R1911 vss.n1140 vss.n1127 2.46896
R1912 vss.n1154 vss.n1153 2.46896
R1913 vss.n52 vss.n51 2.46896
R1914 vss.n46 vss.n10 2.46896
R1915 vss.n44 vss.n43 2.46896
R1916 vss.n39 vss.n38 2.46896
R1917 vss.n36 vss.n35 2.46896
R1918 vss.n31 vss.n30 2.46896
R1919 vss.n28 vss.n27 2.46896
R1920 vss.n23 vss.n22 2.46896
R1921 vss.n20 vss.n19 2.46896
R1922 vss.n1150 vss.n1149 2.46896
R1923 vss.n1147 vss.n1144 2.46896
R1924 vss.n1160 vss.n1159 2.46896
R1925 vss.n1142 vss.n1139 2.46896
R1926 vss.n1168 vss.n1167 2.46896
R1927 vss.n1173 vss.n1172 2.46896
R1928 vss.n1137 vss.n1136 2.46896
R1929 vss.n1132 vss.n58 2.46896
R1930 vss.n1680 vss.n1679 2.46896
R1931 vss.n1683 vss.n1682 2.46896
R1932 vss.n722 vss.n694 2.46896
R1933 vss.n1042 vss.n1041 2.4353
R1934 vss.n1043 vss.n1042 2.4353
R1935 vss.n1546 vss.n1545 2.43106
R1936 vss.n1387 vss.n1386 2.34587
R1937 vss.n1564 vss.t2 2.29252
R1938 vss.n1289 vss.n1288 2.24677
R1939 vss.n318 vss.n246 2.21884
R1940 vss.n1592 vss.n1591 2.21684
R1941 vss.n317 vss.n245 2.18241
R1942 vss.n1339 vss.n417 2.09769
R1943 vss.n1348 vss.n417 2.09769
R1944 vss.n649 vss.n545 2.09769
R1945 vss.n640 vss.n545 2.09769
R1946 vss.n845 vss.n844 2.09769
R1947 vss.n1083 vss.n436 2.09769
R1948 vss.n1605 vss.n206 2.0756
R1949 vss.n155 vss.n148 2.05118
R1950 vss.n168 vss.n153 2.05118
R1951 vss.n168 vss.n154 2.05118
R1952 vss.n161 vss.n148 2.05118
R1953 vss.n169 vss.n168 2.05118
R1954 vss.n156 vss.n148 2.05118
R1955 vss.n170 vss.n148 2.05118
R1956 vss.n1485 vss.n1484 2.05118
R1957 vss.n372 vss.n355 2.05118
R1958 vss.n377 vss.n355 2.05118
R1959 vss.n1484 vss.n358 2.05118
R1960 vss.n382 vss.n355 2.05118
R1961 vss.n1484 vss.n359 2.05118
R1962 vss.n1484 vss.n360 2.05118
R1963 vss.n826 vss.n671 2.03729
R1964 vss.n825 vss.n674 2.03729
R1965 vss.n826 vss.n670 2.03729
R1966 vss.n825 vss.n675 2.03729
R1967 vss.n826 vss.n669 2.03729
R1968 vss.n825 vss.n823 2.03729
R1969 vss.n826 vss.n668 2.03729
R1970 vss.n1306 vss.n1303 2.02871
R1971 vss.n1233 vss.n1232 1.93435
R1972 vss.n1232 vss.n527 1.93435
R1973 vss.n1292 vss.n1291 1.85424
R1974 vss.n236 vss.n235 1.78186
R1975 vss.n1290 vss.n1289 1.76262
R1976 vss.n323 vss.n204 1.76161
R1977 vss.n1548 vss.n1547 1.76161
R1978 vss.n650 vss.n633 1.73826
R1979 vss.n843 vss.n635 1.73826
R1980 vss.n636 vss.n634 1.73826
R1981 vss.n1098 vss.n1097 1.73826
R1982 vss.n1099 vss.n1075 1.73826
R1983 vss.n1103 vss.n1072 1.73826
R1984 vss.n1350 vss.n1349 1.73826
R1985 vss.n1355 vss.n447 1.73826
R1986 vss.n1358 vss.n445 1.73826
R1987 vss.n1290 vss.n466 1.72019
R1988 vss.n1601 vss.n220 1.71592
R1989 vss.n1589 vss.n222 1.71592
R1990 vss.n1585 vss.n230 1.71592
R1991 vss.n1549 vss.n323 1.67978
R1992 vss.n237 vss.n236 1.67978
R1993 vss.n1547 vss.n1546 1.67978
R1994 vss.n236 vss.n228 1.67978
R1995 vss.n1291 vss.n505 1.67438
R1996 vss.n1232 vss.n1231 1.63433
R1997 vss.n1212 vss.n56 1.62307
R1998 vss.n1498 vss.n322 1.39647
R1999 vss.n1042 vss.n1040 1.38385
R2000 vss.n943 vss.n942 1.36702
R2001 vss.n944 vss.n943 1.36702
R2002 vss.n1018 vss.n937 1.36702
R2003 vss.n1018 vss.n936 1.36702
R2004 vss.n979 vss.n978 1.36702
R2005 vss.n980 vss.n979 1.36702
R2006 vss.n1000 vss.n973 1.36702
R2007 vss.n1000 vss.n972 1.36702
R2008 vss.n1493 vss.n204 1.36702
R2009 vss.n1577 vss.n1575 1.36702
R2010 vss.n1567 vss.n244 1.36702
R2011 vss.n265 vss.n233 1.36702
R2012 vss.n303 vss.n302 1.36702
R2013 vss.n288 vss.n256 1.36702
R2014 vss.n1658 vss.n83 1.36702
R2015 vss.n144 vss.n100 1.36702
R2016 vss.n138 vss.n137 1.36702
R2017 vss.n138 vss.n123 1.36702
R2018 vss.n138 vss.n122 1.36702
R2019 vss.n138 vss.n121 1.36702
R2020 vss.n1364 vss.n401 1.36702
R2021 vss.n1373 vss.n1372 1.36702
R2022 vss.n1117 vss.n1116 1.36702
R2023 vss.n1199 vss.n1198 1.36702
R2024 vss.n1499 vss.n330 1.36702
R2025 vss.n1505 vss.n330 1.36702
R2026 vss.n1496 vss.n330 1.36702
R2027 vss.n1517 vss.n1490 1.36702
R2028 vss.n1406 vss.n1405 1.36702
R2029 vss.n745 vss.n744 1.36702
R2030 vss.n779 vss.n737 1.36702
R2031 vss.n877 vss.n559 1.36702
R2032 vss.n866 vss.n559 1.36702
R2033 vss.n902 vss.n901 1.36702
R2034 vss.n902 vss.n560 1.36702
R2035 vss.n902 vss.n561 1.36702
R2036 vss.n902 vss.n562 1.36702
R2037 vss.n902 vss.n563 1.36702
R2038 vss.n902 vss.n564 1.36702
R2039 vss.n902 vss.n565 1.36702
R2040 vss.n903 vss.n902 1.36702
R2041 vss.n610 vss.n572 1.36702
R2042 vss.n610 vss.n573 1.36702
R2043 vss.n610 vss.n583 1.36702
R2044 vss.n610 vss.n584 1.36702
R2045 vss.n610 vss.n585 1.36702
R2046 vss.n610 vss.n586 1.36702
R2047 vss.n610 vss.n587 1.36702
R2048 vss.n610 vss.n609 1.36702
R2049 vss.n707 vss.n625 1.36702
R2050 vss.n1272 vss.n6 1.36702
R2051 vss.n1265 vss.n6 1.36702
R2052 vss.n1263 vss.n6 1.36702
R2053 vss.n1257 vss.n6 1.36702
R2054 vss.n1255 vss.n6 1.36702
R2055 vss.n1249 vss.n6 1.36702
R2056 vss.n1247 vss.n6 1.36702
R2057 vss.n1241 vss.n6 1.36702
R2058 vss.n1239 vss.n6 1.36702
R2059 vss.n1307 vss.n1306 1.36702
R2060 vss.n1306 vss.n473 1.36702
R2061 vss.n1125 vss.n529 1.36702
R2062 vss.n1188 vss.n75 1.36702
R2063 vss.n1179 vss.n1178 1.36702
R2064 vss.n1179 vss.n1127 1.36702
R2065 vss.n1155 vss.n1154 1.36702
R2066 vss.n51 vss.n5 1.36702
R2067 vss.n10 vss.n5 1.36702
R2068 vss.n44 vss.n5 1.36702
R2069 vss.n38 vss.n5 1.36702
R2070 vss.n36 vss.n5 1.36702
R2071 vss.n30 vss.n5 1.36702
R2072 vss.n28 vss.n5 1.36702
R2073 vss.n22 vss.n5 1.36702
R2074 vss.n20 vss.n5 1.36702
R2075 vss.n1149 vss.n56 1.36702
R2076 vss.n1147 vss.n56 1.36702
R2077 vss.n1159 vss.n56 1.36702
R2078 vss.n1142 vss.n56 1.36702
R2079 vss.n1167 vss.n56 1.36702
R2080 vss.n1172 vss.n56 1.36702
R2081 vss.n1137 vss.n56 1.36702
R2082 vss.n1132 vss.n56 1.36702
R2083 vss.n1679 vss.n56 1.36702
R2084 vss.n1682 vss.n56 1.36702
R2085 vss.n722 vss.n721 1.36702
R2086 vss.n641 vss.n624 1.34665
R2087 vss.n1088 vss.n1087 1.34665
R2088 vss.n1341 vss.n1340 1.34665
R2089 vss.n138 vss.n112 1.29223
R2090 vss.n504 vss.n466 1.27538
R2091 vss.n493 vss.n466 1.27538
R2092 vss.n491 vss.n466 1.27538
R2093 vss.n485 vss.n466 1.27538
R2094 vss.n1312 vss.n466 1.27538
R2095 vss.n1315 vss.n466 1.27538
R2096 vss.n1278 vss.n466 1.27538
R2097 vss.n1281 vss.n466 1.27538
R2098 vss.n1617 vss.n1616 1.21742
R2099 vss.n1606 vss.n218 1.21742
R2100 vss.n1600 vss.n223 1.21742
R2101 vss.n310 vss.n309 1.21742
R2102 vss.n1055 vss.n1054 1.21742
R2103 vss.n1036 vss.n0 1.1995
R2104 vss.n1692 vss.n0 1.1365
R2105 vss.n1302 vss.n479 1.13204
R2106 vss.n1388 vss.n441 1.13204
R2107 vss.n1381 vss.n409 1.13204
R2108 vss.n1436 vss.n409 1.13204
R2109 vss.n1449 vss.n369 1.13204
R2110 vss.n1477 vss.n369 1.13204
R2111 vss.n1473 vss.n388 1.13204
R2112 vss.n1543 vss.n326 1.13204
R2113 vss.n676 vss.n668 1.12841
R2114 vss.n823 vss.n822 1.12841
R2115 vss.n819 vss.n669 1.12841
R2116 vss.n817 vss.n675 1.12841
R2117 vss.n815 vss.n670 1.12841
R2118 vss.n813 vss.n674 1.12841
R2119 vss.n672 vss.n671 1.12841
R2120 vss.n813 vss.n671 1.12841
R2121 vss.n815 vss.n674 1.12841
R2122 vss.n817 vss.n670 1.12841
R2123 vss.n819 vss.n675 1.12841
R2124 vss.n822 vss.n669 1.12841
R2125 vss.n823 vss.n676 1.12841
R2126 vss.n824 vss.n668 1.12841
R2127 vss.n1605 vss.n220 1.10722
R2128 vss.n1601 vss.n222 1.10722
R2129 vss.n1589 vss.n230 1.10722
R2130 vss.n1585 vss.n232 1.10722
R2131 vss.n167 vss.n155 1.10063
R2132 vss.n164 vss.n153 1.10063
R2133 vss.n161 vss.n160 1.10063
R2134 vss.n160 vss.n154 1.10063
R2135 vss.n156 vss.n152 1.10063
R2136 vss.n169 vss.n152 1.10063
R2137 vss.n170 vss.n97 1.10063
R2138 vss.n1486 vss.n1485 1.10063
R2139 vss.n372 vss.n356 1.10063
R2140 vss.n376 vss.n358 1.10063
R2141 vss.n377 vss.n376 1.10063
R2142 vss.n381 vss.n359 1.10063
R2143 vss.n382 vss.n381 1.10063
R2144 vss.n385 vss.n360 1.10063
R2145 vss.n164 vss.n155 1.10063
R2146 vss.n162 vss.n153 1.10063
R2147 vss.n162 vss.n161 1.10063
R2148 vss.n157 vss.n154 1.10063
R2149 vss.n157 vss.n156 1.10063
R2150 vss.n171 vss.n169 1.10063
R2151 vss.n171 vss.n170 1.10063
R2152 vss.n1485 vss.n356 1.10063
R2153 vss.n373 vss.n372 1.10063
R2154 vss.n373 vss.n358 1.10063
R2155 vss.n378 vss.n377 1.10063
R2156 vss.n378 vss.n359 1.10063
R2157 vss.n383 vss.n382 1.10063
R2158 vss.n383 vss.n360 1.10063
R2159 vss.n1473 vss.n370 1.09876
R2160 vss.n1036 vss.n1035 1.0945
R2161 vss.n846 vss.n845 1.00762
R2162 vss.n641 vss.n640 1.00762
R2163 vss.n649 vss.n648 1.00762
R2164 vss.n1083 vss.n1082 1.00762
R2165 vss.n1348 vss.n1347 1.00762
R2166 vss.n1339 vss.n1338 1.00762
R2167 vss.n1340 vss.n1339 1.00762
R2168 vss.n1349 vss.n1348 1.00762
R2169 vss.n640 vss.n639 1.00762
R2170 vss.n650 vss.n649 1.00762
R2171 vss.n845 vss.n632 1.00762
R2172 vss.n1084 vss.n1083 1.00762
R2173 vss.n646 vss.n624 0.93057
R2174 vss.n647 vss.n646 0.93057
R2175 vss.n1080 vss.n73 0.93057
R2176 vss.n1087 vss.n1080 0.93057
R2177 vss.n1342 vss.n449 0.93057
R2178 vss.n1342 vss.n1341 0.93057
R2179 vss.n1613 vss.n212 0.919358
R2180 vss.n1298 vss.n479 0.832513
R2181 vss.n1297 vss.n437 0.832513
R2182 vss.n1392 vss.n438 0.832513
R2183 vss.n1040 vss.n6 0.811783
R2184 vss.n1393 vss.n436 0.811783
R2185 vss.n388 vss.n348 0.788139
R2186 vss.n1522 vss.n345 0.788139
R2187 vss.n1528 vss.n346 0.788139
R2188 vss.n795 vss.n794 0.784993
R2189 vss.n307 vss.n306 0.784504
R2190 vss.n1595 vss.n1592 0.769314
R2191 vss.n1592 vss.n227 0.769314
R2192 vss.n635 vss.n633 0.759241
R2193 vss.n843 vss.n636 0.759241
R2194 vss.n838 vss.n634 0.759241
R2195 vss.n1099 vss.n1098 0.759241
R2196 vss.n1103 vss.n1075 0.759241
R2197 vss.n1106 vss.n1072 0.759241
R2198 vss.n1350 vss.n447 0.759241
R2199 vss.n1355 vss.n445 0.759241
R2200 vss.n1359 vss.n1358 0.759241
R2201 vss.n997 vss 0.752
R2202 vss.n1440 vss.n408 0.721578
R2203 vss.n1445 vss.n397 0.721578
R2204 vss.n1449 vss.n395 0.721578
R2205 vss.n1122 vss.n1069 0.6815
R2206 vss.n1215 vss.n506 0.679605
R2207 vss.n1563 vss.n1562 0.672217
R2208 vss.n798 vss 0.661349
R2209 vss.n1511 vss.n1510 0.645237
R2210 vss.n1385 vss.n443 0.621736
R2211 vss.n731 vss.n730 0.619705
R2212 vss.n846 vss.n631 0.587913
R2213 vss.n1082 vss.n79 0.587913
R2214 vss.n1334 vss.n456 0.587913
R2215 vss.n1563 vss.n237 0.583833
R2216 vss.n1206 vss.n1069 0.5675
R2217 vss.n1038 vss.n1037 0.55402
R2218 vss.n1544 vss.n1543 0.544082
R2219 vss.n639 vss.n632 0.538962
R2220 vss.n1085 vss.n1084 0.538962
R2221 vss.n1338 vss.n453 0.538962
R2222 vss.n1386 vss.n1385 0.511252
R2223 vss.n1386 vss.n441 0.511252
R2224 vss.n1381 vss.n443 0.510801
R2225 vss vss.n542 0.478625
R2226 vss.n1564 vss.n226 0.475206
R2227 vss.n774 vss.n735 0.470735
R2228 vss.n1013 vss.n1012 0.450745
R2229 vss.n1031 vss.n1030 0.450745
R2230 vss.n1034 vss.n1033 0.444875
R2231 vss.n1037 vss.n541 0.434812
R2232 vss.n752 vss.n748 0.426816
R2233 vss.n1215 vss.n476 0.422053
R2234 vss.n1545 vss.n1544 0.422053
R2235 vss.n1436 vss.n408 0.41096
R2236 vss.n1440 vss.n397 0.41096
R2237 vss.n1445 vss.n395 0.41096
R2238 vss.n1211 vss.n529 0.406142
R2239 vss.n1286 vss.n509 0.406142
R2240 vss.t76 vss.n466 0.406142
R2241 vss.n1666 vss.t72 0.406142
R2242 vss.n1399 vss.n426 0.406142
R2243 vss.t37 vss.n435 0.406142
R2244 vss.n686 vss 0.396648
R2245 vss.n299 vss.n298 0.386553
R2246 vss.n313 vss 0.38075
R2247 vss.n1664 vss.n1663 0.379017
R2248 vss.n1323 vss.n1322 0.379017
R2249 vss.n850 vss.n849 0.379017
R2250 vss.n1120 vss.n1119 0.376364
R2251 vss.n756 vss.n740 0.349842
R2252 vss.n1639 vss.n107 0.346289
R2253 vss.n766 vss.n765 0.346289
R2254 vss.n1522 vss.n348 0.344399
R2255 vss.n1528 vss.n345 0.344399
R2256 vss.n346 vss.n326 0.344399
R2257 vss.n916 vss.n914 0.338
R2258 vss.n1685 vss.n1684 0.338
R2259 vss.n1686 vss.n54 0.338
R2260 vss.n1284 vss.n1283 0.338
R2261 vss.n1275 vss.n1274 0.338
R2262 vss.n613 vss.n570 0.338
R2263 vss.n899 vss.n614 0.338
R2264 vss vss.n226 0.337094
R2265 vss.n308 vss 0.336026
R2266 vss.n308 vss.n307 0.325763
R2267 vss.n719 vss.n718 0.308395
R2268 vss.n1033 vss 0.307625
R2269 vss.n1185 vss.n1068 0.302237
R2270 vss.n270 vss 0.302
R2271 vss.n1298 vss.n1297 0.300025
R2272 vss.n1392 vss.n437 0.300025
R2273 vss.n1388 vss.n438 0.300025
R2274 vss.n300 vss.n262 0.29236
R2275 vss.n989 vss.n987 0.283526
R2276 vss.n983 vss.n982 0.283526
R2277 vss.n953 vss.n951 0.283526
R2278 vss.n947 vss.n946 0.283526
R2279 vss.n1123 vss.n1121 0.282239
R2280 vss vss.n995 0.279745
R2281 vss vss.n959 0.279745
R2282 vss.n997 vss 0.255875
R2283 vss.n1015 vss 0.255875
R2284 vss vss.n1034 0.255875
R2285 vss.n1121 vss.n1067 0.231731
R2286 vss.n918 vss.n917 0.228708
R2287 vss.n711 vss.n700 0.216049
R2288 vss.n293 vss.n292 0.216026
R2289 vss.n294 vss.n293 0.216026
R2290 vss.n1193 vss.n1192 0.201292
R2291 vss.n285 vss.n264 0.201292
R2292 vss vss.n726 0.193682
R2293 vss.n728 vss.n686 0.182778
R2294 vss.n1518 vss.n1517 0.181328
R2295 vss vss.n996 0.179375
R2296 vss vss.n1014 0.179375
R2297 vss vss.n1032 0.179375
R2298 vss.n1228 vss.n531 0.174427
R2299 vss.n704 vss.n703 0.172625
R2300 vss.n831 vss.n830 0.171026
R2301 vss.n848 vss.n629 0.171026
R2302 vss.n1662 vss.n1661 0.171026
R2303 vss.n106 vss.n105 0.171026
R2304 vss.n1641 vss.n106 0.171026
R2305 vss.n313 vss.n252 0.171026
R2306 vss.n293 vss.n263 0.171026
R2307 vss.n455 vss.n454 0.171026
R2308 vss.n1488 vss.n352 0.171026
R2309 vss.n1489 vss.n1488 0.171026
R2310 vss.n830 vss.n829 0.171026
R2311 vss.n790 vss.n789 0.171026
R2312 vss.n1581 vss.n1580 0.168686
R2313 vss.n1039 vss.n1038 0.166654
R2314 vss.n752 vss.n751 0.164429
R2315 vss.n751 vss.n750 0.164429
R2316 vss.n728 vss.n727 0.163682
R2317 vss.n1598 vss.n1597 0.163106
R2318 vss.n1676 vss.n1675 0.161799
R2319 vss.n1319 vss.n1318 0.161799
R2320 vss.n894 vss.n893 0.161799
R2321 vss.n1014 vss.n1013 0.16025
R2322 vss.n1032 vss.n1031 0.16025
R2323 vss.n1206 vss.n2 0.147897
R2324 vss.n648 vss.n647 0.147353
R2325 vss.n1077 vss.n73 0.147353
R2326 vss.n1347 vss.n449 0.147353
R2327 vss.n191 vss.n190 0.146252
R2328 vss.n1194 vss.n1193 0.145456
R2329 vss.n1195 vss.n87 0.145456
R2330 vss.n730 vss.n684 0.144974
R2331 vss.n729 vss.n685 0.144974
R2332 vss.n1412 vss.n1411 0.144974
R2333 vss.n307 vss.n258 0.144974
R2334 vss.n1059 vss.n1056 0.144974
R2335 vss.n1015 vss 0.143375
R2336 vss.n725 vss.n691 0.143064
R2337 vss.n725 vss.n724 0.142605
R2338 vss.n998 vss.n997 0.142605
R2339 vss.n1006 vss.n1005 0.142605
R2340 vss.n1016 vss.n1015 0.142605
R2341 vss.n1034 vss.n543 0.142605
R2342 vss.n1024 vss.n1023 0.142605
R2343 vss.n1208 vss.n1067 0.141731
R2344 vss.n729 vss.n728 0.141409
R2345 vss.n90 vss.n87 0.140677
R2346 vss vss.n731 0.134375
R2347 vss.n306 vss 0.134375
R2348 vss.n1572 vss.n1571 0.131835
R2349 vss.n1632 vss.n116 0.130763
R2350 vss.n1236 vss.n1235 0.130656
R2351 vss.n1571 vss.n1570 0.127559
R2352 vss.n705 vss.n704 0.127211
R2353 vss.n1193 vss.n1118 0.127211
R2354 vss.n1656 vss.n86 0.127211
R2355 vss.n1654 vss.n87 0.127211
R2356 vss.n182 vss.n181 0.127211
R2357 vss.n192 vss.n191 0.127211
R2358 vss.n277 vss.n264 0.127211
R2359 vss.n1631 vss.n117 0.127211
R2360 vss.n1623 vss.n1622 0.127211
R2361 vss.n1558 vss.n243 0.127211
R2362 vss.n1559 vss.n1558 0.127211
R2363 vss.n995 vss.n994 0.126026
R2364 vss.n1012 vss.n961 0.126026
R2365 vss.n959 vss.n958 0.126026
R2366 vss.n1030 vss.n925 0.126026
R2367 vss.n1691 vss.n1 0.122474
R2368 vss.n191 vss.n142 0.122358
R2369 vss.n1622 vss.n199 0.122358
R2370 vss.n1622 vss.n1621 0.122358
R2371 vss.n280 vss.n264 0.122358
R2372 vss.n269 vss.n251 0.121833
R2373 vss.n314 vss.n313 0.121833
R2374 vss.n313 vss.n312 0.121833
R2375 vss.n724 vss.n692 0.121289
R2376 vss.n719 vss.n692 0.121289
R2377 vss.n718 vss.n717 0.121289
R2378 vss.n701 vss.n700 0.121289
R2379 vss.n705 vss.n701 0.121289
R2380 vss.n994 vss.n993 0.121289
R2381 vss.n993 vss.n990 0.121289
R2382 vss.n990 vss.n989 0.121289
R2383 vss.n984 vss.n983 0.121289
R2384 vss.n986 vss.n984 0.121289
R2385 vss.n987 vss.n986 0.121289
R2386 vss.n976 vss.n961 0.121289
R2387 vss.n976 vss.n974 0.121289
R2388 vss.n982 vss.n974 0.121289
R2389 vss.n958 vss.n957 0.121289
R2390 vss.n957 vss.n954 0.121289
R2391 vss.n954 vss.n953 0.121289
R2392 vss.n948 vss.n947 0.121289
R2393 vss.n950 vss.n948 0.121289
R2394 vss.n951 vss.n950 0.121289
R2395 vss.n940 vss.n925 0.121289
R2396 vss.n940 vss.n938 0.121289
R2397 vss.n946 vss.n938 0.121289
R2398 vss.n832 vss.n831 0.121289
R2399 vss.n832 vss.n629 0.121289
R2400 vss.n917 vss.n916 0.121289
R2401 vss.n581 vss.n580 0.121289
R2402 vss.n580 vss.n579 0.121289
R2403 vss.n579 vss.n576 0.121289
R2404 vss.n576 vss.n575 0.121289
R2405 vss.n575 vss.n553 0.121289
R2406 vss.n913 vss.n553 0.121289
R2407 vss.n914 vss.n913 0.121289
R2408 vss.n1186 vss.n1185 0.121289
R2409 vss.n1186 vss.n1118 0.121289
R2410 vss.n1684 vss.n55 0.121289
R2411 vss.n57 vss.n55 0.121289
R2412 vss.n1677 vss.n57 0.121289
R2413 vss.n1686 vss.n1685 0.121289
R2414 vss.n54 vss.n53 0.121289
R2415 vss.n53 vss.n9 0.121289
R2416 vss.n48 vss.n9 0.121289
R2417 vss.n48 vss.n47 0.121289
R2418 vss.n47 vss.n11 0.121289
R2419 vss.n42 vss.n11 0.121289
R2420 vss.n42 vss.n41 0.121289
R2421 vss.n41 vss.n40 0.121289
R2422 vss.n40 vss.n13 0.121289
R2423 vss.n34 vss.n13 0.121289
R2424 vss.n34 vss.n33 0.121289
R2425 vss.n33 vss.n32 0.121289
R2426 vss.n32 vss.n15 0.121289
R2427 vss.n26 vss.n15 0.121289
R2428 vss.n26 vss.n25 0.121289
R2429 vss.n25 vss.n24 0.121289
R2430 vss.n24 vss.n17 0.121289
R2431 vss.n18 vss.n17 0.121289
R2432 vss.n18 vss.n1 0.121289
R2433 vss.n1183 vss.n1182 0.121289
R2434 vss.n1192 vss.n1183 0.121289
R2435 vss.n1661 vss.n78 0.121289
R2436 vss.n105 vss.n78 0.121289
R2437 vss.n1641 vss.n1640 0.121289
R2438 vss.n1640 vss.n1639 0.121289
R2439 vss.n125 vss.n107 0.121289
R2440 vss.n128 vss.n125 0.121289
R2441 vss.n129 vss.n128 0.121289
R2442 vss.n132 vss.n129 0.121289
R2443 vss.n133 vss.n132 0.121289
R2444 vss.n134 vss.n133 0.121289
R2445 vss.n134 vss.n116 0.121289
R2446 vss.n1656 vss.n1655 0.121289
R2447 vss.n1655 vss.n1654 0.121289
R2448 vss.n181 vss.n145 0.121289
R2449 vss.n192 vss.n145 0.121289
R2450 vss.n263 vss.n252 0.121289
R2451 vss.n286 vss.n285 0.121289
R2452 vss.n292 vss.n286 0.121289
R2453 vss.n295 vss.n294 0.121289
R2454 vss.n298 vss.n295 0.121289
R2455 vss.n300 vss.n299 0.121289
R2456 vss.n276 vss.n266 0.121289
R2457 vss.n277 vss.n276 0.121289
R2458 vss.n1624 vss.n117 0.121289
R2459 vss.n1624 vss.n1623 0.121289
R2460 vss.n454 vss.n404 0.121289
R2461 vss.n404 vss.n352 0.121289
R2462 vss.n1519 vss.n1489 0.121289
R2463 vss.n1519 vss.n1518 0.121289
R2464 vss.n1580 vss.n1579 0.121289
R2465 vss.n1579 vss.n243 0.121289
R2466 vss.n1573 vss.n1559 0.121289
R2467 vss.n1573 vss.n1572 0.121289
R2468 vss.n1283 vss.n1276 0.121289
R2469 vss.n1277 vss.n1276 0.121289
R2470 vss.n1277 vss.n463 0.121289
R2471 vss.n1284 vss.n1275 0.121289
R2472 vss.n1274 vss.n513 0.121289
R2473 vss.n1269 vss.n513 0.121289
R2474 vss.n1269 vss.n1268 0.121289
R2475 vss.n1268 vss.n1267 0.121289
R2476 vss.n1267 vss.n515 0.121289
R2477 vss.n1261 vss.n515 0.121289
R2478 vss.n1261 vss.n1260 0.121289
R2479 vss.n1260 vss.n1259 0.121289
R2480 vss.n1259 vss.n517 0.121289
R2481 vss.n1253 vss.n517 0.121289
R2482 vss.n1253 vss.n1252 0.121289
R2483 vss.n1252 vss.n1251 0.121289
R2484 vss.n1251 vss.n519 0.121289
R2485 vss.n1245 vss.n519 0.121289
R2486 vss.n1245 vss.n1244 0.121289
R2487 vss.n1244 vss.n1243 0.121289
R2488 vss.n1243 vss.n521 0.121289
R2489 vss.n1237 vss.n521 0.121289
R2490 vss.n1237 vss.n1236 0.121289
R2491 vss.n590 vss.n570 0.121289
R2492 vss.n607 vss.n590 0.121289
R2493 vss.n607 vss.n606 0.121289
R2494 vss.n606 vss.n605 0.121289
R2495 vss.n605 vss.n602 0.121289
R2496 vss.n602 vss.n601 0.121289
R2497 vss.n601 vss.n598 0.121289
R2498 vss.n598 vss.n597 0.121289
R2499 vss.n597 vss.n594 0.121289
R2500 vss.n594 vss.n593 0.121289
R2501 vss.n614 vss.n613 0.121289
R2502 vss.n899 vss.n898 0.121289
R2503 vss.n898 vss.n897 0.121289
R2504 vss.n897 vss.n896 0.121289
R2505 vss.n765 vss.n664 0.121289
R2506 vss.n829 vss.n664 0.121289
R2507 vss.n747 vss.n740 0.121289
R2508 vss.n748 vss.n747 0.121289
R2509 vss.n757 vss.n756 0.121289
R2510 vss.n790 vss.n757 0.121289
R2511 vss.n767 vss.n766 0.121289
R2512 vss.n767 vss.n759 0.121289
R2513 vss.n788 vss.n759 0.121289
R2514 vss.n1207 vss.n1068 0.120962
R2515 vss.n717 vss.n697 0.119987
R2516 vss.n1674 vss.n60 0.119721
R2517 vss.n1664 vss.n60 0.119721
R2518 vss.n1324 vss.n1320 0.119721
R2519 vss.n1324 vss.n1323 0.119721
R2520 vss.n850 vss.n616 0.119721
R2521 vss.n892 vss.n616 0.119721
R2522 vss.n1039 vss.n531 0.118192
R2523 vss.n703 vss.n697 0.11525
R2524 vss.n1235 vss.n1234 0.112224
R2525 vss.n1229 vss.n1228 0.112224
R2526 vss.n763 vss.n762 0.104479
R2527 vss.n1123 vss.n1122 0.100283
R2528 vss.n730 vss.n729 0.0982273
R2529 vss.n726 vss.n725 0.0973182
R2530 vss.n593 vss.n541 0.0928684
R2531 vss.n1552 vss.n322 0.0925455
R2532 vss.n1631 vss.n1630 0.0923
R2533 vss.n1570 vss.n1560 0.0905
R2534 vss.n1565 vss.n1560 0.0905
R2535 vss.n1045 vss.n1038 0.0857632
R2536 vss.n1677 vss.n1676 0.0839545
R2537 vss.n1318 vss.n463 0.0839545
R2538 vss.n896 vss.n894 0.0839545
R2539 vss.n1196 vss.n1194 0.0817389
R2540 vss.n1196 vss.n1195 0.0817389
R2541 vss.n146 vss.n91 0.0817389
R2542 vss.n189 vss.n146 0.0817389
R2543 vss.n190 vss.n189 0.0817389
R2544 vss.n197 vss.n142 0.0817389
R2545 vss.n198 vss.n197 0.0817389
R2546 vss.n199 vss.n198 0.0817389
R2547 vss.n1621 vss.n200 0.0817389
R2548 vss.n279 vss.n200 0.0817389
R2549 vss.n280 vss.n279 0.0817389
R2550 vss.n1234 vss.n524 0.0796379
R2551 vss.n1229 vss.n524 0.0796379
R2552 vss.n777 vss.n772 0.076587
R2553 vss.n1632 vss.n1631 0.0736303
R2554 vss.n235 vss.n234 0.0719375
R2555 vss.n271 vss.n270 0.0695
R2556 vss.n315 vss.n251 0.0685
R2557 vss.n315 vss.n314 0.0685
R2558 vss.n312 vss.n253 0.0685
R2559 vss.n262 vss.n253 0.0685
R2560 vss.n1691 vss.n1690 0.068186
R2561 vss.n1235 vss.n523 0.0667727
R2562 vss.n1122 vss.n1120 0.0664166
R2563 vss.n1228 vss.n1227 0.0663636
R2564 vss.n1597 vss.n225 0.0641432
R2565 vss.n1558 vss.n1557 0.0630909
R2566 vss.n1630 vss.n118 0.0617
R2567 vss.n268 vss.n118 0.0617
R2568 vss.n271 vss.n268 0.0617
R2569 vss.n1516 vss.n1515 0.061494
R2570 vss.n1663 vss.n1662 0.0598265
R2571 vss.n1322 vss.n455 0.0598265
R2572 vss.n849 vss.n848 0.0598265
R2573 vss.n713 vss.n691 0.0597258
R2574 vss.n713 vss.n712 0.0597258
R2575 vss.n712 vss.n711 0.0597258
R2576 vss.n643 vss.n623 0.0596781
R2577 vss.n888 vss.n887 0.0596781
R2578 vss.n1670 vss.n69 0.0596781
R2579 vss.n488 vss.n459 0.0596781
R2580 vss.n1091 vss.n72 0.0572123
R2581 vss.n1345 vss.n450 0.0572123
R2582 vss.n1302 vss.n476 0.0559675
R2583 vss.n727 vss 0.0545909
R2584 vss vss.n1596 0.0545
R2585 vss.n830 vss.n663 0.0542097
R2586 vss.n995 vss.n969 0.0525435
R2587 vss.n959 vss.n933 0.0525435
R2588 vss.n166 vss.n106 0.0525312
R2589 vss.n1488 vss.n1487 0.0525312
R2590 vss.n659 vss.n658 0.0524302
R2591 vss vss.n734 0.0518423
R2592 vss.n1571 vss.n231 0.0503024
R2593 vss.n269 vss.n266 0.0502368
R2594 vss.n811 vss.n806 0.0500277
R2595 vss.n811 vss.n810 0.0500277
R2596 vss.n1046 vss.n1045 0.0488158
R2597 vss.n1061 vss.n1046 0.0488158
R2598 vss.n1061 vss.n1060 0.0488158
R2599 vss.n1058 vss.n424 0.0488158
R2600 vss.n1401 vss.n424 0.0488158
R2601 vss.n1402 vss.n1401 0.0488158
R2602 vss.n1403 vss.n421 0.0488158
R2603 vss.n1408 vss.n421 0.0488158
R2604 vss.n1409 vss.n1408 0.0488158
R2605 vss.n1418 vss.n1417 0.0488158
R2606 vss.n1417 vss.n1416 0.0488158
R2607 vss.n1416 vss.n1413 0.0488158
R2608 vss.n1453 vss.n391 0.0488158
R2609 vss.n1454 vss.n1453 0.0488158
R2610 vss.n1455 vss.n1454 0.0488158
R2611 vss.n1458 vss.n1455 0.0488158
R2612 vss.n1457 vss.n1456 0.0488158
R2613 vss.n1456 vss.n334 0.0488158
R2614 vss.n334 vss.n331 0.0488158
R2615 vss.n1539 vss.n332 0.0488158
R2616 vss.n332 vss.n225 0.0488158
R2617 vss.n749 vss.n735 0.0487143
R2618 vss.n1059 vss.n1058 0.0473947
R2619 vss vss.n1692 0.0435
R2620 vss.n855 vss.n623 0.0424178
R2621 vss.n888 vss.n855 0.0424178
R2622 vss.n1670 vss.n1669 0.0424178
R2623 vss.n1669 vss.n1668 0.0424178
R2624 vss.n1327 vss.n459 0.0424178
R2625 vss.n1328 vss.n1327 0.0424178
R2626 vss.n1134 vss.n59 0.0422273
R2627 vss.n1170 vss.n1138 0.0422273
R2628 vss.n1170 vss.n1169 0.0422273
R2629 vss.n1165 vss.n1164 0.0422273
R2630 vss.n1552 vss.n319 0.0422273
R2631 vss.n1556 vss.n319 0.0422273
R2632 vss.n1557 vss.n1556 0.0422273
R2633 vss.n1317 vss.n464 0.0422273
R2634 vss.n487 vss.n470 0.0422273
R2635 vss.n489 vss.n487 0.0422273
R2636 vss.n495 vss.n483 0.0422273
R2637 vss.n1218 vss.n1217 0.0422273
R2638 vss.n1608 vss.n216 0.0422273
R2639 vss.n859 vss.n615 0.0422273
R2640 vss.n872 vss.n869 0.0422273
R2641 vss.n873 vss.n872 0.0422273
R2642 vss.n886 vss.n883 0.0422273
R2643 vss.n906 vss.n905 0.0422273
R2644 vss.n908 vss.n906 0.0422273
R2645 vss.n908 vss.n907 0.0422273
R2646 vss.n1157 vss.n1156 0.0416619
R2647 vss.n1295 vss.n1294 0.0414091
R2648 vss.n812 vss.n811 0.0404194
R2649 vss.n1004 vss.n969 0.040413
R2650 vss.n1022 vss.n933 0.040413
R2651 vss.n184 vss.n173 0.0391719
R2652 vss.n1475 vss.n386 0.0391719
R2653 vss vss.n659 0.0389394
R2654 vss.n1690 vss.n2 0.0384339
R2655 vss.n677 vss.n663 0.0375161
R2656 vss.n821 vss.n677 0.0375161
R2657 vss.n821 vss.n820 0.0375161
R2658 vss.n820 vss.n818 0.0375161
R2659 vss.n818 vss.n816 0.0375161
R2660 vss.n816 vss.n814 0.0375161
R2661 vss.n814 vss.n812 0.0375161
R2662 vss vss.n1457 0.0374474
R2663 vss.n1012 vss 0.0368913
R2664 vss.n1030 vss 0.0368913
R2665 vss.n166 vss.n165 0.0363594
R2666 vss.n165 vss.n163 0.0363594
R2667 vss.n163 vss.n159 0.0363594
R2668 vss.n159 vss.n158 0.0363594
R2669 vss.n158 vss.n151 0.0363594
R2670 vss.n172 vss.n151 0.0363594
R2671 vss.n173 vss.n172 0.0363594
R2672 vss.n1487 vss.n353 0.0363594
R2673 vss.n374 vss.n353 0.0363594
R2674 vss.n375 vss.n374 0.0363594
R2675 vss.n379 vss.n375 0.0363594
R2676 vss.n380 vss.n379 0.0363594
R2677 vss.n384 vss.n380 0.0363594
R2678 vss.n386 vss.n384 0.0363594
R2679 vss.n1165 vss.n69 0.0360909
R2680 vss.n488 vss.n483 0.0360909
R2681 vss.n887 vss.n886 0.0360909
R2682 vss.n1413 vss.n1412 0.0360263
R2683 vss.n1108 vss.n1107 0.0351154
R2684 vss.n1383 vss.n1360 0.0351154
R2685 vss.n839 vss.n659 0.0351154
R2686 vss.n1410 vss.n1409 0.0341316
R2687 vss.n1477 vss.n370 0.0337805
R2688 vss.n1005 vss.n968 0.0337609
R2689 vss.n1023 vss.n932 0.0337609
R2690 vss.n1081 vss.n77 0.0325979
R2691 vss.n1089 vss.n1086 0.0325979
R2692 vss.n1092 vss.n1089 0.0325979
R2693 vss.n1090 vss.n1078 0.0325979
R2694 vss.n1336 vss.n1335 0.0325979
R2695 vss.n1337 vss.n451 0.0325979
R2696 vss.n1344 vss.n451 0.0325979
R2697 vss.n1346 vss.n448 0.0325979
R2698 vss.n847 vss.n630 0.0325979
R2699 vss.n642 vss.n638 0.0325979
R2700 vss.n644 vss.n642 0.0325979
R2701 vss.n651 vss.n637 0.0325979
R2702 vss.n1121 vss.n1069 0.0323462
R2703 vss.n1210 vss.n508 0.032
R2704 vss.n1224 vss.n532 0.0315909
R2705 vss.n1223 vss.n535 0.0315909
R2706 vss.n1052 vss.n538 0.0315909
R2707 vss.n1051 vss.n1050 0.0315909
R2708 vss.n1049 vss.n1048 0.0315909
R2709 vss.n1397 vss.n430 0.0315909
R2710 vss.n1396 vss.n431 0.0315909
R2711 vss.n1370 vss.n434 0.0315909
R2712 vss.n1369 vss.n1368 0.0315909
R2713 vss.n1375 vss.n1366 0.0315909
R2714 vss.n1377 vss.n1376 0.0315909
R2715 vss.n1378 vss.n416 0.0315909
R2716 vss.n415 vss.n412 0.0315909
R2717 vss.n1433 vss.n1432 0.0315909
R2718 vss.n1429 vss.n413 0.0315909
R2719 vss.n1428 vss.n1427 0.0315909
R2720 vss.n1426 vss.n1425 0.0315909
R2721 vss.n1481 vss.n364 0.0315909
R2722 vss.n1480 vss.n365 0.0315909
R2723 vss.n1469 vss.n1463 0.0315909
R2724 vss.n1468 vss.n1466 0.0315909
R2725 vss.n1465 vss.n1464 0.0315909
R2726 vss.n1533 vss.n339 0.0315909
R2727 vss.n1532 vss.n342 0.0315909
R2728 vss.n341 vss.n340 0.0315909
R2729 vss.n1611 vss.n215 0.0315909
R2730 vss.n1610 vss.n1609 0.0315909
R2731 vss.n1604 vss.n207 0.0310309
R2732 vss.n1540 vss.n1539 0.0293947
R2733 vss.n1134 vss.n1133 0.0291364
R2734 vss.n1176 vss.n1130 0.0291364
R2735 vss.n1175 vss.n1131 0.0291364
R2736 vss.n1304 vss.n464 0.0291364
R2737 vss.n469 vss.n467 0.0291364
R2738 vss.n1310 vss.n1309 0.0291364
R2739 vss.n860 vss.n859 0.0291364
R2740 vss.n864 vss.n863 0.0291364
R2741 vss.n868 vss.n856 0.0291364
R2742 vss.n1515 vss.n1492 0.0281506
R2743 vss.n1492 vss.n242 0.0281506
R2744 vss.n1581 vss.n242 0.0281506
R2745 vss.n654 vss.n552 0.0271119
R2746 vss.n918 vss.n552 0.0266818
R2747 vss.n1206 vss.n1205 0.0264129
R2748 vss vss.n1402 0.0260789
R2749 vss.n270 vss.n269 0.0258333
R2750 vss.n1164 vss.n1163 0.0254545
R2751 vss.n1162 vss.n1141 0.0254545
R2752 vss.n1145 vss.n1143 0.0254545
R2753 vss.n498 vss.n495 0.0254545
R2754 vss.n501 vss.n499 0.0254545
R2755 vss.n502 vss.n481 0.0254545
R2756 vss.n883 vss.n874 0.0254545
R2757 vss.n880 vss.n879 0.0254545
R2758 vss.n875 vss.n557 0.0254545
R2759 vss.n1091 vss.n1090 0.0247308
R2760 vss.n1346 vss.n1345 0.0247308
R2761 vss.n643 vss.n637 0.0247308
R2762 vss.n1516 vss.n1491 0.0242273
R2763 vss.n968 vss.n962 0.023587
R2764 vss.n932 vss.n926 0.023587
R2765 vss.n183 vss.n182 0.0232801
R2766 vss.n1403 vss 0.0232368
R2767 vss.n1078 vss.n1076 0.0228427
R2768 vss.n1101 vss.n1100 0.0228427
R2769 vss.n1102 vss.n1071 0.0228427
R2770 vss.n1351 vss.n448 0.0228427
R2771 vss.n1354 vss.n1352 0.0228427
R2772 vss.n1353 vss.n444 0.0228427
R2773 vss.n652 vss.n651 0.0228427
R2774 vss.n842 vss.n653 0.0228427
R2775 vss.n841 vss.n840 0.0228427
R2776 vss.n1501 vss.n322 0.0225909
R2777 vss.n1603 vss.n1602 0.0225553
R2778 vss.n1588 vss.n221 0.0225553
R2779 vss.n1587 vss.n1586 0.0225553
R2780 vss.n1508 vss.n1507 0.0221818
R2781 vss.n1503 vss.n1495 0.0221818
R2782 vss.n1502 vss.n1501 0.0221818
R2783 vss.n1208 vss.n1207 0.0212692
R2784 vss.n789 vss.n758 0.0209545
R2785 vss.n734 vss.n678 0.0206745
R2786 vss.n581 vss.n541 0.0206316
R2787 vss.n1508 vss.n1491 0.0205455
R2788 vss.n1507 vss.n1495 0.0205455
R2789 vss.n1503 vss.n1502 0.0205455
R2790 vss.n1207 vss.n1206 0.0202191
R2791 vss.n1517 vss.n1516 0.0200181
R2792 vss.n1540 vss.n331 0.0199211
R2793 vss.n806 vss.n805 0.0193501
R2794 vss.n810 vss.n807 0.0193501
R2795 vss.n807 vss.n661 0.0193501
R2796 vss.n657 vss.n656 0.0193501
R2797 vss.n656 vss.n654 0.0193501
R2798 vss.n1596 vss.n226 0.0190625
R2799 vss.n1597 vss 0.0176913
R2800 vss.n1011 vss.n962 0.0173261
R2801 vss.n1029 vss.n926 0.0173261
R2802 vss.n1163 vss.n1162 0.0172727
R2803 vss.n1143 vss.n1141 0.0172727
R2804 vss.n1157 vss.n1145 0.0172727
R2805 vss.n499 vss.n498 0.0172727
R2806 vss.n502 vss.n501 0.0172727
R2807 vss.n1294 vss.n481 0.0172727
R2808 vss.n880 vss.n874 0.0172727
R2809 vss.n879 vss.n875 0.0172727
R2810 vss.n905 vss.n557 0.0172727
R2811 vss.n789 vss.n788 0.0171646
R2812 vss.n324 vss.n322 0.0168636
R2813 vss.n805 vss.n678 0.0164061
R2814 vss vss.n1011 0.0161522
R2815 vss vss.n1029 0.0161522
R2816 vss.n907 vss.n552 0.0160455
R2817 vss.n782 vss.n773 0.0155852
R2818 vss.n781 vss.n778 0.0155852
R2819 vss.n776 vss.n774 0.0155852
R2820 vss.n1418 vss.n1410 0.0151842
R2821 vss.n661 vss 0.0150996
R2822 vss.n1384 vss.n440 0.0150483
R2823 vss.n1382 vss.n1361 0.0150483
R2824 vss.n1448 vss.n371 0.0150483
R2825 vss.n1476 vss.n371 0.0150483
R2826 vss.n1474 vss.n387 0.0150483
R2827 vss.n1525 vss.n327 0.0150483
R2828 vss.n327 vss.n208 0.0150483
R2829 vss.n1301 vss.n1300 0.0150483
R2830 vss.n1389 vss.n440 0.0150483
R2831 vss.n1604 vss.n1603 0.0147292
R2832 vss.n1602 vss.n221 0.0147292
R2833 vss.n1588 vss.n1587 0.0147292
R2834 vss.n1586 vss.n231 0.0147292
R2835 vss.n1475 vss.n1474 0.0146204
R2836 vss.n1133 vss.n1130 0.0135909
R2837 vss.n1176 vss.n1175 0.0135909
R2838 vss.n1138 vss.n1131 0.0135909
R2839 vss.n1304 vss.n467 0.0135909
R2840 vss.n1310 vss.n469 0.0135909
R2841 vss.n1309 vss.n470 0.0135909
R2842 vss.n863 vss.n860 0.0135909
R2843 vss.n864 vss.n856 0.0135909
R2844 vss.n869 vss.n868 0.0135909
R2845 vss.n794 vss.n735 0.0134262
R2846 vss.n1152 vss.n1146 0.0133933
R2847 vss.n1146 vss.n1070 0.0133933
R2848 vss.n1412 vss.n391 0.0132895
R2849 vss.n1114 vss.n1112 0.0131971
R2850 vss.n185 vss.n95 0.0131971
R2851 vss.n1634 vss.n1633 0.0131971
R2852 vss.n1114 vss 0.0130726
R2853 vss.n94 vss.n86 0.0129481
R2854 vss.n1218 vss.n505 0.0128745
R2855 vss.n1204 vss.n1108 0.0125747
R2856 vss.n1458 vss 0.0118684
R2857 vss.n773 vss.n758 0.0114943
R2858 vss.n782 vss.n781 0.0114943
R2859 vss.n778 vss.n776 0.0114943
R2860 vss.n1301 vss.n1295 0.0114826
R2861 vss.n185 vss.n184 0.0113299
R2862 vss.n1300 vss.n1299 0.0111973
R2863 vss.n1296 vss.n439 0.0111973
R2864 vss.n1391 vss.n1390 0.0111973
R2865 vss.n1227 vss.n532 0.0111364
R2866 vss.n1224 vss.n1223 0.0111364
R2867 vss.n538 vss.n535 0.0111364
R2868 vss.n1052 vss.n1051 0.0111364
R2869 vss.n1050 vss.n1049 0.0111364
R2870 vss.n1048 vss.n430 0.0111364
R2871 vss.n1397 vss.n1396 0.0111364
R2872 vss.n434 vss.n431 0.0111364
R2873 vss.n1370 vss.n1369 0.0111364
R2874 vss.n1368 vss.n1366 0.0111364
R2875 vss.n1376 vss.n1375 0.0111364
R2876 vss.n1378 vss.n1377 0.0111364
R2877 vss.n416 vss.n415 0.0111364
R2878 vss.n1433 vss.n412 0.0111364
R2879 vss.n1432 vss.n413 0.0111364
R2880 vss.n1429 vss.n1428 0.0111364
R2881 vss.n1427 vss.n1426 0.0111364
R2882 vss.n1425 vss.n364 0.0111364
R2883 vss.n1481 vss.n1480 0.0111364
R2884 vss.n1463 vss.n365 0.0111364
R2885 vss.n1469 vss.n1468 0.0111364
R2886 vss.n1466 vss.n1465 0.0111364
R2887 vss.n1464 vss.n339 0.0111364
R2888 vss.n1533 vss.n1532 0.0111364
R2889 vss.n342 vss.n341 0.0111364
R2890 vss.n340 vss.n215 0.0111364
R2891 vss.n1611 vss.n1610 0.0111364
R2892 vss.n1609 vss.n1608 0.0111364
R2893 vss.n1088 vss.n1079 0.0108879
R2894 vss.n1648 vss.n94 0.010832
R2895 vss.n1647 vss.n95 0.010832
R2896 vss.n1548 vss.n324 0.0107694
R2897 vss.n1210 vss.n523 0.0107273
R2898 vss.n1217 vss.n508 0.0107273
R2899 vss.n387 vss.n347 0.0106268
R2900 vss.n1524 vss.n1523 0.0106268
R2901 vss.n1527 vss.n1526 0.0106268
R2902 vss.n234 vss.n226 0.010625
R2903 vss vss.n1113 0.010334
R2904 vss.n176 vss.n99 0.010334
R2905 vss.n175 vss.n174 0.010334
R2906 vss.n1634 vss.n115 0.010334
R2907 vss.n1100 vss.n1076 0.0102552
R2908 vss.n1102 vss.n1101 0.0102552
R2909 vss.n1107 vss.n1071 0.0102552
R2910 vss.n1352 vss.n1351 0.0102552
R2911 vss.n1354 vss.n1353 0.0102552
R2912 vss.n1360 vss.n444 0.0102552
R2913 vss.n653 vss.n652 0.0102552
R2914 vss.n842 vss.n841 0.0102552
R2915 vss.n840 vss.n839 0.0102552
R2916 vss.n750 vss.n749 0.0101429
R2917 vss.n1439 vss.n1438 0.009771
R2918 vss.n1446 vss.n396 0.009771
R2919 vss.n1448 vss.n1447 0.009771
R2920 vss.n182 vss.n99 0.00971162
R2921 vss.n1361 vss 0.00905784
R2922 vss.n1155 vss.n1152 0.0088427
R2923 vss.n1384 vss.n1383 0.00848732
R2924 vss.n1092 vss.n1091 0.00836713
R2925 vss.n1345 vss.n1344 0.00836713
R2926 vss.n644 vss.n643 0.00836713
R2927 vss.n1662 vss.n77 0.00805245
R2928 vss.n1335 vss.n455 0.00805245
R2929 vss.n848 vss.n847 0.00805245
R2930 vss.n1182 vss.n1119 0.00760526
R2931 vss.n1675 vss.n1674 0.00751299
R2932 vss.n1320 vss.n1319 0.00751299
R2933 vss.n893 vss.n892 0.00751299
R2934 vss.n1086 vss.n1081 0.00742308
R2935 vss.n1337 vss.n1336 0.00742308
R2936 vss.n638 vss.n630 0.00742308
R2937 vss.n1205 vss.n1070 0.00732584
R2938 vss.n505 vss.n480 0.00720365
R2939 vss.n1005 vss.n1004 0.00715217
R2940 vss.n1023 vss.n1022 0.00715217
R2941 vss.n1383 vss.n1382 0.00706101
R2942 vss.n1169 vss.n69 0.00663636
R2943 vss.n489 vss.n488 0.00663636
R2944 vss.n887 vss.n873 0.00663636
R2945 vss.n1437 vss 0.00649049
R2946 vss.n1205 vss.n1204 0.00622614
R2947 vss.n91 vss.n90 0.00607522
R2948 vss.n235 vss.n216 0.00581818
R2949 vss.n1565 vss.n1564 0.00579412
R2950 vss.n1438 vss.n1437 0.00577734
R2951 vss.n1439 vss.n396 0.00577734
R2952 vss.n1447 vss.n1446 0.00577734
R2953 vss.n1156 vss.n1155 0.00505056
R2954 vss.n1523 vss.n347 0.00492155
R2955 vss.n1527 vss.n1524 0.00492155
R2956 vss.n1526 vss.n1525 0.00492155
R2957 vss.n1299 vss.n1296 0.00435103
R2958 vss.n1391 vss.n439 0.00435103
R2959 vss.n1390 vss.n1389 0.00435103
R2960 vss.n1295 vss.n480 0.00406577
R2961 vss.n176 vss.n175 0.00336307
R2962 vss.n174 vss.n115 0.00336307
R2963 vss.n324 vss.n208 0.00320998
R2964 vss.n1668 vss.n72 0.00296575
R2965 vss.n1328 vss.n450 0.00296575
R2966 vss.n1676 vss.n59 0.00295455
R2967 vss.n1318 vss.n1317 0.00295455
R2968 vss.n894 vss.n615 0.00295455
R2969 vss.n1648 vss.n1647 0.00286515
R2970 vss.n184 vss.n183 0.00236722
R2971 vss.n1548 vss.n207 0.00206894
R2972 vss.n735 vss 0.00194966
R2973 vss.n1060 vss.n1059 0.00192105
R2974 vss.n658 vss.n657 0.00160883
R2975 vss.n1112 vss.n1108 0.00112241
R2976 vss.n1476 vss.n1475 0.000927892
R2977 vss.n1113 vss.n86 0.000748963
R2978 vss.n1633 vss.n1632 0.000624481
R2979 vdd.t45 vdd.t62 933.037
R2980 vdd.t62 vdd.t64 834.822
R2981 vdd.t25 vdd.t11 715.827
R2982 vdd.t6 vdd.t20 594.059
R2983 vdd.n166 vdd.t29 501.8
R2984 vdd.n103 vdd.t10 501.8
R2985 vdd.t10 vdd 489.991
R2986 vdd.n169 vdd.t29 489.502
R2987 vdd.n167 vdd.t25 489.219
R2988 vdd.n33 vdd.t27 489.219
R2989 vdd.n63 vdd.t3 476.993
R2990 vdd.t11 vdd.n166 476.62
R2991 vdd.t20 vdd.n103 476.62
R2992 vdd.t27 vdd.n32 336.332
R2993 vdd.n57 vdd.n53 330.935
R2994 vdd.t68 vdd.n58 311.151
R2995 vdd.t3 vdd.t21 306.656
R2996 vdd.n45 vdd.n42 277.878
R2997 vdd.n39 vdd.t58 266.188
R2998 vdd.n105 vdd.n104 256.137
R2999 vdd.n30 vdd.t0 250.899
R3000 vdd.n36 vdd.t0 244.75
R3001 vdd.n47 vdd.t51 238.31
R3002 vdd.n50 vdd.t66 238.31
R3003 vdd.t14 vdd.n51 238.31
R3004 vdd.n62 vdd.t52 238.31
R3005 vdd.t60 vdd.n40 215.827
R3006 vdd.t47 vdd.t60 215.827
R3007 vdd.t16 vdd.t54 201.44
R3008 vdd.t51 vdd.n46 197.843
R3009 vdd.t18 vdd.t23 191.548
R3010 vdd.n41 vdd.t12 178.958
R3011 vdd.n52 vdd.t5 178.059
R3012 vdd.t56 vdd.n45 160.072
R3013 vdd.n46 vdd.t48 160.072
R3014 vdd.t50 vdd.t47 142.087
R3015 vdd.t44 vdd.t8 131.296
R3016 vdd.t1 vdd.t68 126.799
R3017 vdd.n61 vdd.n59 126.799
R3018 vdd.t52 vdd.n61 124.102
R3019 vdd.n104 vdd.t6 117.007
R3020 vdd.n59 vdd.t1 111.511
R3021 vdd.n32 vdd.t44 107.014
R3022 vdd.t8 vdd.n30 107.014
R3023 vdd.t54 vdd.t14 102.519
R3024 vdd.n51 vdd.n50 90.8278
R3025 vdd.t48 vdd.t56 78.2379
R3026 vdd.t21 vdd.n62 69.2451
R3027 vdd.n12 vdd.n11 62.0058
R3028 vdd.n146 vdd.n145 62.0058
R3029 vdd.n94 vdd.n93 62.0058
R3030 vdd.n104 vdd.t45 60.2684
R3031 vdd.n53 vdd.n52 60.2523
R3032 vdd.t12 vdd.t50 59.353
R3033 vdd.n3 vdd.n2 54.711
R3034 vdd.n135 vdd.n134 54.711
R3035 vdd.n125 vdd.n88 54.711
R3036 vdd.n109 vdd.n101 54.5452
R3037 vdd.n110 vdd.n109 54.5452
R3038 vdd.t5 vdd.t16 53.9573
R3039 vdd.n42 vdd.n41 53.0581
R3040 vdd.n111 vdd.n110 48.3037
R3041 vdd.t23 vdd.n57 46.7631
R3042 vdd.n58 vdd.t18 46.7631
R3043 vdd.n7 vdd.n6 44.4321
R3044 vdd.n21 vdd.n7 44.4321
R3045 vdd.n139 vdd.n138 44.4321
R3046 vdd.n155 vdd.n139 44.4321
R3047 vdd.n123 vdd.n89 44.4321
R3048 vdd.n124 vdd.n123 44.4321
R3049 vdd.n14 vdd.n13 44.1177
R3050 vdd.n148 vdd.n147 44.1177
R3051 vdd.n117 vdd.n116 41.0086
R3052 vdd.n14 vdd.n5 31.6537
R3053 vdd.n148 vdd.n137 31.6537
R3054 vdd.n118 vdd.n117 31.6537
R3055 vdd.n13 vdd.n12 29.9841
R3056 vdd.n147 vdd.n146 29.9841
R3057 vdd.n115 vdd.n93 29.9841
R3058 vdd.n6 vdd.n2 29.5043
R3059 vdd.n138 vdd.n134 29.5043
R3060 vdd.n125 vdd.n124 29.5043
R3061 vdd.n101 vdd.n92 28.5602
R3062 vdd.n161 vdd.t40 26.892
R3063 vdd.n141 vdd.t34 24.3938
R3064 vdd.n23 vdd.n22 23.3768
R3065 vdd.n157 vdd.n156 23.3768
R3066 vdd.n91 vdd.n87 23.3768
R3067 vdd.n40 vdd.n39 22.4825
R3068 vdd.n170 vdd.n169 20.3863
R3069 vdd.n84 vdd.n36 20.2319
R3070 vdd.n11 vdd.n3 19.8952
R3071 vdd.n145 vdd.n135 19.8952
R3072 vdd.n94 vdd.n88 19.8952
R3073 vdd vdd.n141 19.301
R3074 vdd.n165 vdd.n164 19.1102
R3075 vdd.n84 vdd 18.6524
R3076 vdd.n29 vdd.n28 18.5371
R3077 vdd.n162 vdd.n161 18.4336
R3078 vdd.n28 vdd.n27 18.3436
R3079 vdd.n164 vdd.n163 18.3436
R3080 vdd.n130 vdd.n129 18.3436
R3081 vdd.n131 vdd.n130 18.3166
R3082 vdd.n27 vdd.t37 13.1071
R3083 vdd.n163 vdd.t39 13.1071
R3084 vdd.n141 vdd.t35 13.1071
R3085 vdd.n129 vdd.t33 13.1071
R3086 vdd.n168 vdd.n166 12.8823
R3087 vdd.n103 vdd.n102 12.8823
R3088 vdd.n64 vdd.n62 12.8823
R3089 vdd.n67 vdd.n59 12.8823
R3090 vdd.n71 vdd.n53 12.8823
R3091 vdd.n80 vdd.n41 12.8823
R3092 vdd.n72 vdd.n52 12.8823
R3093 vdd.n79 vdd.n42 12.8823
R3094 vdd vdd.n47 12.8823
R3095 vdd.n35 vdd.n30 12.8823
R3096 vdd.n40 vdd.n38 12.6005
R3097 vdd.n46 vdd.n44 12.6005
R3098 vdd.n50 vdd.n48 12.6005
R3099 vdd.n58 vdd.n55 12.6005
R3100 vdd.n61 vdd.n60 12.6005
R3101 vdd.n39 vdd.n37 12.6005
R3102 vdd.n45 vdd.n43 12.6005
R3103 vdd.n51 vdd.n49 12.6005
R3104 vdd.n57 vdd.n54 12.6005
R3105 vdd.n32 vdd.n31 12.6005
R3106 vdd.n161 vdd.t41 10.8823
R3107 vdd.n22 vdd.n4 10.8334
R3108 vdd.n156 vdd.n136 10.8334
R3109 vdd.n95 vdd.n91 10.8334
R3110 vdd.n10 vdd.n4 9.75782
R3111 vdd.n24 vdd.n23 9.75782
R3112 vdd.n144 vdd.n136 9.75782
R3113 vdd.n158 vdd.n157 9.75782
R3114 vdd.n126 vdd.n87 9.75782
R3115 vdd.n96 vdd.n95 9.75782
R3116 vdd vdd.t53 9.21665
R3117 vdd.n16 vdd.t43 8.94208
R3118 vdd.n17 vdd.t42 8.94208
R3119 vdd.n150 vdd.t31 8.94208
R3120 vdd.n151 vdd.t30 8.94208
R3121 vdd.n100 vdd.t63 8.94208
R3122 vdd.n121 vdd.t65 8.94208
R3123 vdd.n63 vdd.t4 8.42234
R3124 vdd.n65 vdd.t22 8.42234
R3125 vdd.n73 vdd.t17 8.42234
R3126 vdd.n74 vdd.t55 8.42234
R3127 vdd.n81 vdd.t13 8.42234
R3128 vdd.n167 vdd.t26 8.31339
R3129 vdd.n105 vdd.t7 8.31339
R3130 vdd.n54 vdd.t19 8.31339
R3131 vdd.n49 vdd.t15 8.31339
R3132 vdd.n43 vdd.t49 8.31339
R3133 vdd.n37 vdd.t61 8.31339
R3134 vdd.n31 vdd.t9 8.31339
R3135 vdd.n33 vdd.t28 8.31339
R3136 vdd.n60 vdd.t2 8.30475
R3137 vdd.n55 vdd.t24 8.30475
R3138 vdd.n48 vdd.t67 8.30475
R3139 vdd.n44 vdd.t57 8.30475
R3140 vdd.n38 vdd.t59 8.30475
R3141 vdd.n56 vdd.t69 8.1405
R3142 vdd.n23 vdd.n3 6.79787
R3143 vdd.n157 vdd.n135 6.79787
R3144 vdd.n88 vdd.n87 6.79787
R3145 vdd.n111 vdd.n92 4.97256
R3146 vdd.n22 vdd.n21 3.64787
R3147 vdd.n156 vdd.n155 3.64787
R3148 vdd.n91 vdd.n89 3.64787
R3149 vdd.n113 vdd.t46 3.52948
R3150 vdd.n116 vdd.n115 3.23339
R3151 vdd.n11 vdd.n4 3.1505
R3152 vdd.n145 vdd.n136 3.1505
R3153 vdd.n95 vdd.n94 3.1505
R3154 vdd.n27 vdd.t36 2.24244
R3155 vdd.n163 vdd.t38 2.24244
R3156 vdd.n129 vdd.t32 2.24244
R3157 vdd.n13 vdd.n8 2.1005
R3158 vdd.n21 vdd.n20 2.1005
R3159 vdd.n20 vdd.n5 2.1005
R3160 vdd.n6 vdd.n0 2.1005
R3161 vdd.n147 vdd.n140 2.1005
R3162 vdd.n155 vdd.n154 2.1005
R3163 vdd.n154 vdd.n137 2.1005
R3164 vdd.n138 vdd.n132 2.1005
R3165 vdd.n115 vdd.n114 2.1005
R3166 vdd.n124 vdd.n85 2.1005
R3167 vdd.n119 vdd.n118 2.1005
R3168 vdd.n119 vdd.n89 2.1005
R3169 vdd.t66 vdd.n47 1.79906
R3170 vdd.n22 vdd.n5 1.69074
R3171 vdd.n156 vdd.n137 1.69074
R3172 vdd.n118 vdd.n91 1.69074
R3173 vdd.n15 vdd.n14 1.5755
R3174 vdd.n18 vdd.n7 1.5755
R3175 vdd.n25 vdd.n24 1.5755
R3176 vdd.n10 vdd.n9 1.5755
R3177 vdd.n149 vdd.n148 1.5755
R3178 vdd.n152 vdd.n139 1.5755
R3179 vdd.n144 vdd.n143 1.5755
R3180 vdd.n159 vdd.n158 1.5755
R3181 vdd.n106 vdd.n101 1.5755
R3182 vdd.n110 vdd.n99 1.5755
R3183 vdd.n123 vdd.n122 1.5755
R3184 vdd.n117 vdd.n90 1.5755
R3185 vdd.n127 vdd.n126 1.5755
R3186 vdd.n97 vdd.n96 1.5755
R3187 vdd.n12 vdd.n10 1.46026
R3188 vdd.n24 vdd.n2 1.46026
R3189 vdd.n146 vdd.n144 1.46026
R3190 vdd.n158 vdd.n134 1.46026
R3191 vdd.n126 vdd.n125 1.46026
R3192 vdd.n96 vdd.n93 1.46026
R3193 vdd.n131 vdd.n84 1.286
R3194 vdd vdd.n29 1.2385
R3195 vdd.n165 vdd.n131 1.207
R3196 vdd.n112 vdd.n111 1.05197
R3197 vdd.n109 vdd.n108 1.0505
R3198 vdd.n168 vdd.n167 0.942415
R3199 vdd.n108 vdd.n99 0.779711
R3200 vdd.n107 vdd.n102 0.643822
R3201 vdd.n113 vdd.n99 0.622211
R3202 vdd.n15 vdd.n8 0.607567
R3203 vdd.n149 vdd.n140 0.607567
R3204 vdd.n34 vdd.n33 0.567196
R3205 vdd.n142 vdd 0.566593
R3206 vdd.n116 vdd.n92 0.538578
R3207 vdd.n108 vdd.n107 0.512741
R3208 vdd.n28 vdd 0.498918
R3209 vdd.n130 vdd 0.498918
R3210 vdd.n17 vdd.n0 0.48464
R3211 vdd.n151 vdd.n132 0.48464
R3212 vdd.n121 vdd.n85 0.48226
R3213 vdd.n56 vdd 0.395064
R3214 vdd.n9 vdd.n8 0.392291
R3215 vdd vdd.n170 0.3665
R3216 vdd.n169 vdd 0.319524
R3217 vdd.n107 vdd.n105 0.309149
R3218 vdd.n26 vdd.n0 0.285895
R3219 vdd.n142 vdd.n140 0.285895
R3220 vdd.n160 vdd.n132 0.285895
R3221 vdd.n128 vdd.n85 0.285895
R3222 vdd.n19 vdd.n18 0.27928
R3223 vdd.n153 vdd.n152 0.27928
R3224 vdd.n122 vdd.n120 0.275922
R3225 vdd.n120 vdd.n90 0.275922
R3226 vdd.n82 vdd 0.263188
R3227 vdd.n68 vdd.n56 0.26172
R3228 vdd.n70 vdd.n54 0.261195
R3229 vdd.n75 vdd.n49 0.261195
R3230 vdd.n78 vdd.n43 0.261195
R3231 vdd.n83 vdd.n37 0.261195
R3232 vdd.n34 vdd.n31 0.261195
R3233 vdd.n164 vdd 0.247811
R3234 vdd.n36 vdd 0.24575
R3235 vdd.n66 vdd.n60 0.234974
R3236 vdd.n69 vdd.n55 0.234974
R3237 vdd.n76 vdd.n48 0.234974
R3238 vdd.n77 vdd.n44 0.234974
R3239 vdd.n82 vdd.n38 0.234974
R3240 vdd.n35 vdd.n34 0.218188
R3241 vdd.n66 vdd.n65 0.2075
R3242 vdd.n71 vdd.n70 0.205813
R3243 vdd.n79 vdd.n78 0.172625
R3244 vdd.n112 vdd.n100 0.165429
R3245 vdd.n19 vdd.n16 0.156354
R3246 vdd.n153 vdd.n150 0.156354
R3247 vdd vdd.n77 0.150688
R3248 vdd vdd.n76 0.150688
R3249 vdd vdd.n69 0.150688
R3250 vdd.n68 vdd 0.147312
R3251 vdd.n98 vdd.n97 0.138889
R3252 vdd vdd.n74 0.137188
R3253 vdd.n25 vdd.n1 0.136775
R3254 vdd.n9 vdd.n1 0.136775
R3255 vdd.n97 vdd.n86 0.136775
R3256 vdd.n127 vdd.n86 0.136775
R3257 vdd vdd.n83 0.134938
R3258 vdd.n64 vdd 0.132125
R3259 vdd.n74 vdd 0.127063
R3260 vdd.n69 vdd.n68 0.1265
R3261 vdd.n16 vdd.n15 0.123427
R3262 vdd.n18 vdd.n17 0.123427
R3263 vdd.n150 vdd.n149 0.123427
R3264 vdd.n152 vdd.n151 0.123427
R3265 vdd vdd.n102 0.122
R3266 vdd.n122 vdd.n121 0.121946
R3267 vdd.n100 vdd.n90 0.121946
R3268 vdd.n106 vdd.n98 0.117332
R3269 vdd.n120 vdd.n119 0.107
R3270 vdd.n26 vdd.n25 0.106897
R3271 vdd.n128 vdd.n127 0.106897
R3272 vdd.n20 vdd.n19 0.106625
R3273 vdd.n154 vdd.n153 0.106625
R3274 vdd vdd.n26 0.106221
R3275 vdd vdd.n128 0.106221
R3276 vdd.n159 vdd.n133 0.103436
R3277 vdd.n143 vdd.n133 0.103436
R3278 vdd vdd.n81 0.101187
R3279 vdd.n78 vdd 0.101187
R3280 vdd vdd.n73 0.101187
R3281 vdd vdd.n63 0.101187
R3282 vdd.n20 vdd.n1 0.090875
R3283 vdd.n154 vdd.n133 0.090875
R3284 vdd.n119 vdd.n86 0.090875
R3285 vdd.n29 vdd 0.0905
R3286 vdd.n73 vdd.n72 0.082625
R3287 vdd vdd.n162 0.0825588
R3288 vdd.n160 vdd.n159 0.080867
R3289 vdd.n143 vdd.n142 0.080867
R3290 vdd vdd.n168 0.0795244
R3291 vdd vdd.n160 0.0748848
R3292 vdd.n170 vdd.n165 0.072
R3293 vdd vdd.n67 0.071375
R3294 vdd.n67 vdd 0.06125
R3295 vdd vdd.n35 0.06125
R3296 vdd.n76 vdd.n75 0.055625
R3297 vdd.n114 vdd.n113 0.0534573
R3298 vdd.n81 vdd.n80 0.0494375
R3299 vdd.n114 vdd.n98 0.0460488
R3300 vdd.n72 vdd.n71 0.0381875
R3301 vdd.n80 vdd.n79 0.0336875
R3302 vdd.n70 vdd 0.0303125
R3303 vdd.n77 vdd 0.0280625
R3304 vdd.n65 vdd.n64 0.0201875
R3305 vdd vdd.n66 0.0190625
R3306 vdd.n83 vdd.n82 0.01625
R3307 vdd.n75 vdd 0.0156875
R3308 vdd.n107 vdd.n106 0.00329503
R3309 vdd.n162 vdd 0.00201261
R3310 vdd.n113 vdd.n112 0.00187113
R3311 v_rew v_rew.t3 37.2214
R3312 v_rew.n0 v_rew.t0 32.5076
R3313 v_rew.n1 v_rew.t2 28.3362
R3314 v_rew.n2 v_rew.t1 28.3362
R3315 v_rew.n2 v_rew.n1 11.0961
R3316 v_rew.n1 v_rew 5.4005
R3317 v_rew.n0 v_rew 4.71875
R3318 v_rew v_rew.n0 0.104711
R3319 v_rew v_rew.n2 0.102342
R3320 vmem vmem.t0 20.2482
R3321 vmem.n2 vmem.t11 16.4806
R3322 vmem.n2 vmem.n1 14.0833
R3323 vmem.n8 vmem.t10 13.1366
R3324 vmem.n6 vmem.n4 9.716
R3325 vmem.n8 vmem.n7 9.63725
R3326 vmem vmem.t7 9.17794
R3327 vmem vmem.t8 9.14522
R3328 vmem.n6 vmem.n5 9.0005
R3329 vmem.n0 vmem.t6 8.8205
R3330 vmem.n1 vmem.t2 8.8205
R3331 vmem vmem.t4 8.57004
R3332 vmem vmem.t3 8.53506
R3333 vmem.n5 vmem.t5 8.1405
R3334 vmem.n4 vmem.t1 8.1405
R3335 vmem.n3 vmem.n0 5.47925
R3336 vmem.n8 vmem.t9 4.99592
R3337 vmem vmem.n3 4.78962
R3338 vmem.n7 vmem.n6 2.507
R3339 vmem.n7 vmem 2.33487
R3340 vmem.n3 vmem.n2 0.818375
R3341 vmem.n5 vmem 0.427318
R3342 vmem.n0 vmem 0.394944
R3343 vmem.n4 vmem 0.394591
R3344 vmem.n1 vmem 0.323598
R3345 vmem vmem.n8 0.136625
R3346 vin.n0 vin.t4 59.6219
R3347 vin vin.t2 21.3485
R3348 vin.n3 vin.n2 18.652
R3349 vin.n1 vin.n0 18.5261
R3350 vin.n1 vin 12.01
R3351 vin.n3 vin.t1 8.8205
R3352 vin vin.t0 8.54078
R3353 vin vin.n3 0.38923
R3354 vin.n2 vin.t3 0.0455
R3355 vin.n2 vin.n1 0.0305
R3356 vin.n0 vin 0.003875
R3357 phi_fire.n0 phi_fire.t12 41.9396
R3358 phi_fire.n6 phi_fire.t4 41.9396
R3359 phi_fire.n3 phi_fire.t9 39.4319
R3360 phi_fire.n5 phi_fire.t10 37.4396
R3361 phi_fire.n9 phi_fire.t13 37.4396
R3362 phi_fire.n2 phi_fire.t7 34.4873
R3363 phi_fire.n11 phi_fire.t3 33.5205
R3364 phi_fire.n0 phi_fire.t15 32.5076
R3365 phi_fire.n4 phi_fire.t16 32.5076
R3366 phi_fire.n8 phi_fire.t11 32.5076
R3367 phi_fire.n6 phi_fire.t2 32.5076
R3368 phi_fire phi_fire.t6 28.457
R3369 phi_fire.n1 phi_fire.t5 28.3362
R3370 phi_fire.n3 phi_fire.t14 28.3362
R3371 phi_fire.n7 phi_fire.t8 28.3362
R3372 phi_fire.n14 phi_fire 12.9706
R3373 phi_fire.n10 phi_fire.n9 9.9725
R3374 phi_fire phi_fire.n13 9.2525
R3375 phi_fire phi_fire.t0 9.04888
R3376 phi_fire.n12 phi_fire.n11 9.0005
R3377 phi_fire.n14 phi_fire.t1 8.1405
R3378 phi_fire.n12 phi_fire.n5 6.1025
R3379 phi_fire.n10 phi_fire.n7 5.63162
R3380 phi_fire.n2 phi_fire.n1 4.94505
R3381 phi_fire.n5 phi_fire.n4 4.5005
R3382 phi_fire.n9 phi_fire.n8 4.5005
R3383 phi_fire.n13 phi_fire.n12 4.5005
R3384 phi_fire phi_fire.n14 0.332129
R3385 phi_fire.n13 phi_fire.n2 0.321125
R3386 phi_fire.n11 phi_fire.n10 0.255071
R3387 phi_fire phi_fire.n0 0.104711
R3388 phi_fire.n4 phi_fire 0.104711
R3389 phi_fire phi_fire.n6 0.104711
R3390 phi_fire.n1 phi_fire 0.102342
R3391 phi_fire phi_fire.n3 0.102342
R3392 phi_fire.n7 phi_fire 0.102342
R3393 phi_fire.n8 phi_fire 0.0857632
R3394 vout.n0 vout.t2 9.57203
R3395 vout vout.t1 9.21093
R3396 vout.n0 vout.t0 8.1405
R3397 vout.n2 vout.t3 8.1405
R3398 vout.n1 vout.n0 4.84475
R3399 vout.n2 vout.n1 4.5005
R3400 vout.n1 vout 0.856625
R3401 vout vout.n2 0.399071
C0 vmem a_9352_5200# 0.50178f
C1 phi_fire vdd 3.86998f
C2 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.nand$1_0.Z 0.30883f
C3 ota_1stage$2_0.vout a_n872_2246# 0.00619f
C4 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vdd 0.01306f
C5 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.vneg 0.00455f
C6 phaseUpulse_0.vrefrac phaseUpulse_0.phi_2 0.08553f
C7 phaseUpulse_0.monostable_0.nand$1_1.Z v_rew 0.02831f
C8 a_8827_1078# vdd 0.28491f
C9 phaseUpulse_0.conmutator_0.out v_th 0.07509f
C10 a_2328_4757# vdd 0.02704f
C11 vspike phi_fire 0.11476f
C12 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_1 0.36261f
C13 a_2248_2068# phaseUpulse_0.monostable_0.not$1_0.in 0
C14 vspike phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.00386f
C15 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.monostable_0.nand$1_1.Z 0.47242f
C16 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_int 0
C17 a_9352_5200# phi_fire 0.86685f
C18 phaseUpulse_0.vrefrac phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.12269f
C19 v_th phaseUpulse_0.monostable_0.not$1_1.in 0.1654f
C20 vmem v_ref 1.14628f
C21 v_th vdd 0.95711f
C22 phaseUpulse_0.phi_2 v_ref 0.02285f
C23 phaseUpulse_0.conmutator_0.out ota_1stage$2_0.vout 0.00815f
C24 phaseUpulse_0.vrefrac a_2328_4757# 0.24845f
C25 a_2266_6197# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.02959f
C26 v_th v_rew 0.00409f
C27 a_4045_8037# vdd 0.60338f
C28 a_2266_6197# a_2328_4757# 0.37601f
C29 vspike v_th 0.00729f
C30 a_6164_1900# a_6854_3116# 0.47928f
C31 v_ref phi_fire 1.41406f
C32 v_th phaseUpulse_0.monostable_0.not$1_3.in 0.07018f
C33 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp v_ref 0.23381f
C34 ota_1stage$2_0.vout vdd 0.54052f
C35 phaseUpulse_0.vrefrac v_th 0.36994f
C36 a_8811_n132# vin 0.49018f
C37 a_8827_1078# v_ref 0.47663f
C38 a_8190_3623# a_6854_3116# 0.29863f
C39 a_2328_4757# v_ref 0.01863f
C40 ota_1stage$2_0.vout v_rew 0.07589f
C41 a_2521_9609# vdd 1.29114f
C42 a_2266_6197# v_th 0.3674f
C43 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.vspike_down 0.01248f
C44 a_7562_3851# a_6854_3116# 0.39032f
C45 a_8190_3623# a_6164_1900# 0.06628f
C46 vmem conmutator$1_2.out 0.26299f
C47 a_6854_3116# vin 0.21271f
C48 a_3790_4625# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0
C49 ota_1stage$2_0.vout phaseUpulse_0.monostable_0.not$1_3.in 0.01206f
C50 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.monostable_0.not$1_1.in 0.42262f
C51 a_2328_4757# phaseUpulse_0.vspike_down 0
C52 a_7562_3851# a_6164_1900# 0.04031f
C53 phaseUpulse_0.monostable_0.not$1_0.in vdd 0.60484f
C54 v_th v_ref 0.93865f
C55 phaseUpulse_0.monostable_0.nand$1_1.Z a_n1388_602# 0.04857f
C56 a_6164_1900# vin 0.21486f
C57 a_3544_1172# phaseUpulse_0.phi_2 0.01051f
C58 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vneg 0.00125f
C59 a_7562_3851# a_8190_3623# 0.17539f
C60 a_8075_5978# vmem 0.08258f
C61 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vspike_up 0.00609f
C62 a_4045_8037# v_ref 0.00199f
C63 a_8190_3623# vin 0.00184f
C64 a_3790_4625# phaseUpulse_0.vneg 0
C65 conmutator$1_2.out phi_fire 0.61083f
C66 vspike phaseUpulse_0.monostable_0.not$1_0.in 0
C67 v_th phaseUpulse_0.vspike_down 0.27438f
C68 a_8827_1078# conmutator$1_2.out 0.75454f
C69 a_7562_3851# vin 0.11121f
C70 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.vneg 0.00153f
C71 v_th a_1078_602# 0.00317f
C72 phaseUpulse_0.vrefrac phaseUpulse_0.monostable_0.not$1_0.in 0
C73 v_th a_1251_6917# 0.0201f
C74 a_3544_2068# phaseUpulse_0.vneg 0.00155f
C75 a_8075_5978# phi_fire 0.87587f
C76 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_1 0.2402f
C77 phaseUpulse_0.vneg phaseUpulse_0.phi_1 0.37793f
C78 a_2248_2068# phaseUpulse_0.vneg 0.00174f
C79 phaseUpulse_0.vneg phaseUpulse_0.phi_int 0.00786f
C80 ota_1stage$2_0.vout phaseUpulse_0.vspike_down 0
C81 v_th phaseUpulse_0.vspike_up 0.15877f
C82 conmutator$1_0.out vdd 0.41962f
C83 a_3544_2068# phaseUpulse_0.phi_1 0
C84 a_2248_2068# a_3544_2068# 0.00376f
C85 a_3544_2068# phaseUpulse_0.phi_int 0.50615f
C86 phaseUpulse_0.vneg a_n872_2246# 0.02206f
C87 ota_1stage$2_0.vout a_1251_6917# 0
C88 a_2583_8169# vdd 0.06682f
C89 a_2248_2068# phaseUpulse_0.phi_1 0.00836f
C90 a_8811_n132# vdd 0.27677f
C91 phaseUpulse_0.phi_1 phaseUpulse_0.phi_int 0.05163f
C92 a_8190_3623# vout 0.0164f
C93 ota_1stage$2_0.vout a_n1388_602# 0.00427f
C94 a_8075_5978# v_th 0
C95 ota_1stage$2_0.vout phaseUpulse_0.vspike_up 0.58752f
C96 a_6854_3116# vdd 0.06522f
C97 vmem phi_fire 2.73055f
C98 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.phi_2 0.00294f
C99 phaseUpulse_0.monostable_0.not$1_0.in a_1078_602# 0.00381f
C100 vmem a_8827_1078# 0.09883f
C101 a_6164_1900# vdd 0.53169f
C102 phaseUpulse_0.conmutator_0.out phaseUpulse_0.vneg 0.1271f
C103 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn vdd 0.00204f
C104 vspike a_6854_3116# 0.03458f
C105 a_952_2068# v_th 0.01009f
C106 a_8190_3623# vdd 1.10527f
C107 a_3790_4625# vdd 0.57977f
C108 conmutator$1_0.out v_ref 0.05967f
C109 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phi_fire 0.10728f
C110 phaseUpulse_0.conmutator_0.out phaseUpulse_0.phi_1 0.1136f
C111 vspike a_6164_1900# 0.21492f
C112 a_7562_3851# vdd 1.2793f
C113 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.monostable_0.nand$1_0.Z 0.47226f
C114 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.vneg 0
C115 a_8827_1078# phi_fire 0.94674f
C116 phaseUpulse_0.monostable_0.nand$1_0.Z vdd 0.37216f
C117 phaseUpulse_0.vneg vdd 0.84325f
C118 vmem v_th 0.0572f
C119 vdd vin 0.99052f
C120 vspike a_8190_3623# 0.03541f
C121 a_2328_4757# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.05005f
C122 phaseUpulse_0.conmutator_0.out a_n872_2246# 0.83515f
C123 a_3544_2068# vdd 0.27055f
C124 phaseUpulse_0.vrefrac phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0.23309f
C125 phaseUpulse_0.vneg v_rew 0.1251f
C126 a_8190_3623# a_9352_5200# 0.00744f
C127 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_1 0.04237f
C128 vspike a_7562_3851# 0.00374f
C129 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_int 0
C130 phaseUpulse_0.phi_1 vdd 1.6851f
C131 a_2248_2068# vdd 0.27536f
C132 vspike phaseUpulse_0.monostable_0.nand$1_0.Z 0.00176f
C133 a_2266_6197# phaseUpulse_0.refractory_0.ota_1stage$1_0.vn 0.00282f
C134 phaseUpulse_0.vrefrac a_3790_4625# 0.01646f
C135 vspike phaseUpulse_0.vneg 0.0349f
C136 vspike vin 0.18648f
C137 phaseUpulse_0.phi_int vdd 0.70343f
C138 v_th phaseUpulse_0.monostable_0.nand$1_1.Z 0.02529f
C139 a_6854_3116# v_ref 0
C140 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.monostable_0.nand$1_0.Z 0.00483f
C141 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.vneg 0.42522f
C142 vspike a_3544_2068# 0.5989f
C143 v_th phi_fire 0.00717f
C144 phaseUpulse_0.phi_1 v_rew 0.007f
C145 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp v_th 0.00715f
C146 a_n872_2246# vdd 0.75706f
C147 phaseUpulse_0.vrefrac phaseUpulse_0.vneg 0.0665f
C148 a_2266_6197# a_3790_4625# 0.00553f
C149 a_6164_1900# v_ref 0.00178f
C150 vspike phaseUpulse_0.phi_1 0.48921f
C151 vspike a_2248_2068# 0.59888f
C152 a_3544_2068# phaseUpulse_0.vrefrac 0
C153 a_n872_2246# v_rew 0.79579f
C154 a_2328_4757# v_th 0.15887f
C155 vspike phaseUpulse_0.phi_int 0.27454f
C156 a_952_2068# phaseUpulse_0.monostable_0.not$1_0.in 0
C157 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.phi_1 0.00862f
C158 a_8190_3623# v_ref 0.24721f
C159 phaseUpulse_0.vrefrac phaseUpulse_0.phi_1 0.02194f
C160 a_2248_2068# phaseUpulse_0.vrefrac 0.10994f
C161 a_3790_4625# v_ref 0.2647f
C162 phaseUpulse_0.vrefrac phaseUpulse_0.phi_int 0
C163 ota_1stage$2_0.vout phaseUpulse_0.monostable_0.nand$1_1.Z 0.03281f
C164 phaseUpulse_0.monostable_0.not$1_3.in a_n872_2246# 0
C165 conmutator$1_2.out a_8811_n132# 0.0061f
C166 a_7562_3851# v_ref 0
C167 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.vspike_down 0.36026f
C168 vout vdd 0.31925f
C169 phaseUpulse_0.vneg v_ref 0.0771f
C170 phaseUpulse_0.monostable_0.not$1_0.in phaseUpulse_0.phi_2 0.3513f
C171 a_8075_5978# conmutator$1_0.out 0.69525f
C172 v_ref vin 0.0166f
C173 a_3544_2068# v_ref 0.137f
C174 phaseUpulse_0.conmutator_0.out vdd 0.74727f
C175 a_4045_8037# v_th 0
C176 a_6854_3116# conmutator$1_2.out 0.00747f
C177 phaseUpulse_0.conmutator_0.out v_rew 0.75989f
C178 phaseUpulse_0.phi_1 v_ref 0.00326f
C179 a_2248_2068# v_ref 0.01335f
C180 phaseUpulse_0.vneg phaseUpulse_0.vspike_down 0.01362f
C181 phaseUpulse_0.phi_int v_ref 0.23227f
C182 a_9352_5200# vout 0.69632f
C183 a_6164_1900# conmutator$1_2.out 0.03605f
C184 phaseUpulse_0.monostable_0.nand$1_0.Z a_1078_602# 0.04857f
C185 phaseUpulse_0.conmutator_0.out vspike 0.15135f
C186 phaseUpulse_0.monostable_0.not$1_1.in vdd 0.2269f
C187 ota_1stage$2_0.vout v_th 0.0278f
C188 phaseUpulse_0.conmutator_0.out phaseUpulse_0.monostable_0.not$1_3.in 0.00501f
C189 a_8190_3623# conmutator$1_2.out 0.00161f
C190 phaseUpulse_0.conmutator_0.out phaseUpulse_0.vrefrac 0
C191 a_n1388_602# phaseUpulse_0.vneg 0.00381f
C192 v_rew vdd 1.18265f
C193 ota_1stage$2_0.vout a_4045_8037# 0
C194 a_2521_9609# v_th 0.00766f
C195 phaseUpulse_0.phi_1 a_1078_602# 0.00569f
C196 phaseUpulse_0.vneg phaseUpulse_0.vspike_up 0.03807f
C197 a_7562_3851# conmutator$1_2.out 0.00226f
C198 vmem conmutator$1_0.out 0.09392f
C199 vspike phaseUpulse_0.monostable_0.not$1_1.in 0.00276f
C200 vspike vdd 0.89929f
C201 a_2521_9609# a_4045_8037# 0.00553f
C202 conmutator$1_2.out vin 0.79779f
C203 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.monostable_0.not$1_1.in 0.07366f
C204 phaseUpulse_0.monostable_0.not$1_3.in vdd 0.2263f
C205 a_9352_5200# vdd 0.2791f
C206 phaseUpulse_0.vrefrac phaseUpulse_0.monostable_0.not$1_1.in 0
C207 v_ref vout 0.1593f
C208 v_th phaseUpulse_0.monostable_0.not$1_0.in 0.00666f
C209 vmem a_8811_n132# 0.11316f
C210 phaseUpulse_0.vrefrac vdd 0.30981f
C211 a_3544_1172# phaseUpulse_0.vneg 0
C212 phaseUpulse_0.monostable_0.not$1_3.in v_rew 0.0052f
C213 a_3544_2068# a_3544_1172# 0
C214 a_2521_9609# ota_1stage$2_0.vout 0.09327f
C215 conmutator$1_2.out phaseUpulse_0.phi_int 0
C216 a_2266_6197# vdd 1.25241f
C217 conmutator$1_0.out phi_fire 0.55602f
C218 a_n872_2246# phaseUpulse_0.vspike_up 0.08242f
C219 a_3544_1172# phaseUpulse_0.phi_1 0.01f
C220 a_6854_3116# vmem 0.03683f
C221 vspike phaseUpulse_0.vrefrac 0.18182f
C222 a_3544_1172# phaseUpulse_0.phi_int 0.04163f
C223 phi_fire a_8811_n132# 0.54852f
C224 a_6164_1900# vmem 0.1629f
C225 v_ref vdd 0.98376f
C226 a_8827_1078# a_8811_n132# 0
C227 a_952_2068# phaseUpulse_0.monostable_0.nand$1_0.Z 0
C228 a_952_2068# phaseUpulse_0.vneg 0.00415f
C229 a_8190_3623# vmem 1.01491f
C230 a_2266_6197# phaseUpulse_0.vrefrac 0.0563f
C231 a_6854_3116# phi_fire 0.02296f
C232 v_th conmutator$1_0.out 0.05947f
C233 phaseUpulse_0.vspike_down vdd 0.13281f
C234 vspike v_ref 0.2195f
C235 a_7562_3851# vmem 0.01101f
C236 phaseUpulse_0.conmutator_0.out phaseUpulse_0.vspike_up 0.09025f
C237 phaseUpulse_0.monostable_0.not$1_1.in a_1078_602# 0.00369f
C238 a_6164_1900# phi_fire 0.06015f
C239 a_9352_5200# v_ref 0.19585f
C240 phaseUpulse_0.monostable_0.nand$1_0.Z phaseUpulse_0.phi_2 0.00237f
C241 vmem vin 0.35856f
C242 phaseUpulse_0.vneg phaseUpulse_0.phi_2 0.02188f
C243 a_952_2068# phaseUpulse_0.phi_1 0.52142f
C244 a_1078_602# vdd 0.00261f
C245 a_952_2068# a_2248_2068# 0.00376f
C246 v_th a_2583_8169# 0.03955f
C247 a_4045_8037# conmutator$1_0.out 0.09338f
C248 a_1251_6917# vdd 0.00936f
C249 phaseUpulse_0.vrefrac v_ref 0.00382f
C250 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.01318f
C251 a_6164_1900# a_8827_1078# 0.00737f
C252 a_3544_2068# phaseUpulse_0.phi_2 0.0077f
C253 a_8190_3623# phi_fire 0.17771f
C254 a_952_2068# a_n872_2246# 0.00376f
C255 a_4045_8037# a_2583_8169# 0.04633f
C256 a_n1388_602# vdd 0.00261f
C257 a_3790_4625# phi_fire 0.00387f
C258 a_2266_6197# v_ref 0.03181f
C259 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn a_2328_4757# 0.03005f
C260 a_3790_4625# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0.02274f
C261 a_8190_3623# a_8827_1078# 0
C262 phaseUpulse_0.phi_1 phaseUpulse_0.phi_2 0.4489f
C263 a_2248_2068# phaseUpulse_0.phi_2 0.49862f
C264 phaseUpulse_0.vspike_up vdd 0.38521f
C265 a_7562_3851# phi_fire 0.05873f
C266 phaseUpulse_0.vrefrac phaseUpulse_0.vspike_down 0.59606f
C267 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.monostable_0.nand$1_0.Z 0.07835f
C268 phaseUpulse_0.phi_2 phaseUpulse_0.phi_int 0.25422f
C269 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.vneg 0.3112f
C270 a_n1388_602# v_rew 0
C271 conmutator$1_2.out vdd 0.4963f
C272 phaseUpulse_0.vneg phi_fire 0.00133f
C273 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.vneg 0.04823f
C274 a_3790_4625# a_2328_4757# 0.04633f
C275 phi_fire vin 0.28319f
C276 phaseUpulse_0.vspike_up v_rew 0.35339f
C277 ota_1stage$2_0.vout a_2583_8169# 0.21159f
C278 a_2521_9609# conmutator$1_0.out 0.03015f
C279 a_3544_2068# phi_fire 0
C280 phaseUpulse_0.vrefrac a_1251_6917# 0
C281 a_2266_6197# phaseUpulse_0.vspike_down 0.01207f
C282 a_8827_1078# vin 0.00869f
C283 a_3544_1172# vdd 0.05888f
C284 phaseUpulse_0.monostable_0.not$1_3.in a_n1388_602# 0.00369f
C285 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn v_th 0.05102f
C286 phaseUpulse_0.monostable_0.nand$1_1.Z phaseUpulse_0.phi_1 0.00153f
C287 a_2521_9609# a_2583_8169# 0.40678f
C288 phaseUpulse_0.phi_1 phi_fire 0.00103f
C289 a_8075_5978# vdd 0.27975f
C290 vspike conmutator$1_2.out 0.06761f
C291 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.phi_1 0
C292 a_2248_2068# phaseUpulse_0.refractory_0.ota_1stage$1_0.vp 0
C293 phaseUpulse_0.phi_int phi_fire 0.40552f
C294 phaseUpulse_0.monostable_0.not$1_3.in phaseUpulse_0.vspike_up 0
C295 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp phaseUpulse_0.phi_int 0
C296 a_3790_4625# v_th 0.02226f
C297 phaseUpulse_0.vspike_down v_ref 0
C298 phaseUpulse_0.conmutator_0.out a_952_2068# 0.10777f
C299 vspike a_3544_1172# 0.00279f
C300 vmem vout 0.15077f
C301 v_th phaseUpulse_0.monostable_0.nand$1_0.Z 0.17131f
C302 v_th phaseUpulse_0.vneg 0.48308f
C303 v_th vin 0.00917f
C304 a_952_2068# phaseUpulse_0.monostable_0.not$1_1.in 0.0012f
C305 a_952_2068# vdd 0.28111f
C306 v_th phaseUpulse_0.phi_1 0.2582f
C307 a_1251_6917# phaseUpulse_0.vspike_down 0.06482f
C308 phi_fire vout 0.57965f
C309 a_952_2068# v_rew 0.00313f
C310 conmutator$1_2.out v_ref 0.15117f
C311 v_th a_n872_2246# 0
C312 ota_1stage$2_0.vout phaseUpulse_0.vneg 0.20337f
C313 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.phi_2 0.01642f
C314 phaseUpulse_0.conmutator_0.out phaseUpulse_0.monostable_0.nand$1_1.Z 0
C315 vmem vdd 1.21415f
C316 phaseUpulse_0.phi_2 vdd 0.69232f
C317 vspike a_952_2068# 0.55963f
C318 phaseUpulse_0.vspike_up phaseUpulse_0.vspike_down 0.03889f
C319 a_8075_5978# v_ref 0.07879f
C320 a_952_2068# phaseUpulse_0.vrefrac 0.01389f
C321 a_2583_8169# conmutator$1_0.out 0.075f
C322 phaseUpulse_0.vspike_up a_1251_6917# 0.06422f
C323 vspike vmem 0.09386f
C324 phaseUpulse_0.monostable_0.not$1_1.in phaseUpulse_0.monostable_0.nand$1_1.Z 0.00251f
C325 vspike phaseUpulse_0.phi_2 0.27648f
C326 phaseUpulse_0.monostable_0.nand$1_1.Z vdd 0.41173f
C327 v_rew vss 0.82919f
C328 vout vss 0.49719f
C329 vin vss 3.39858f
C330 vdd vss 94.34265f
C331 a_8811_n132# vss 0.20221f
C332 a_1078_602# vss 0.07193f
C333 a_n1388_602# vss 0.07193f
C334 conmutator$1_2.out vss 1.81382f
C335 a_3544_1172# vss 0.00446f
C336 phaseUpulse_0.monostable_0.nand$1_0.Z vss 1.12845f
C337 phaseUpulse_0.monostable_0.nand$1_1.Z vss 1.16177f
C338 a_8827_1078# vss 0.50172f
C339 phaseUpulse_0.monostable_0.not$1_1.in vss 1.45035f
C340 phaseUpulse_0.monostable_0.not$1_0.in vss 0.89494f
C341 phaseUpulse_0.monostable_0.not$1_3.in vss 1.45831f
C342 a_6854_3116# vss 1.2516f
C343 a_6164_1900# vss 2.73439f
C344 a_8190_3623# vss 2.41685f
C345 a_7562_3851# vss 0.56919f
C346 a_3544_2068# vss 0.18952f
C347 a_2248_2068# vss 0.16661f
C348 a_952_2068# vss 0.16613f
C349 vspike vss 2.62702f
C350 phaseUpulse_0.conmutator_0.out vss 0.55274f
C351 phaseUpulse_0.phi_int vss 1.52046f
C352 phaseUpulse_0.phi_2 vss 1.30055f
C353 phaseUpulse_0.phi_1 vss 1.54616f
C354 a_n872_2246# vss 0.52986f
C355 phaseUpulse_0.vneg vss 9.09826f
C356 a_9352_5200# vss 0.49434f
C357 phaseUpulse_0.refractory_0.ota_1stage$1_0.vp vss 3.99233f
C358 a_2328_4757# vss 1.37841f
C359 phaseUpulse_0.refractory_0.ota_1stage$1_0.vn vss 1.5386f
C360 a_3790_4625# vss 1.76476f
C361 phaseUpulse_0.vrefrac vss 1.74013f
C362 a_2266_6197# vss 0.59277f
C363 vmem vss 4.10793f
C364 a_8075_5978# vss 0.956f
C365 phi_fire vss 6.98236f
C366 v_ref vss 5.2017f
C367 phaseUpulse_0.vspike_down vss 2.1272f
C368 a_1251_6917# vss 0.96922f
C369 phaseUpulse_0.vspike_up vss 2.48364f
C370 conmutator$1_0.out vss 3.47422f
C371 a_2583_8169# vss 1.42414f
C372 v_th vss 7.24603f
C373 a_4045_8037# vss 1.87447f
C374 ota_1stage$2_0.vout vss 4.108f
C375 a_2521_9609# vss 0.71365f
C376 phi_fire.t7 vss 0.05811f
C377 phi_fire.t12 vss 0.0516f
C378 phi_fire.t15 vss 0.02985f
C379 phi_fire.n0 vss 0.17293f
C380 phi_fire.t5 vss 0.03833f
C381 phi_fire.n1 vss 0.10909f
C382 phi_fire.n2 vss 0.32578f
C383 phi_fire.t9 vss 0.09582f
C384 phi_fire.t14 vss 0.03833f
C385 phi_fire.n3 vss 0.37206f
C386 phi_fire.t16 vss 0.02985f
C387 phi_fire.n4 vss 0.04111f
C388 phi_fire.t10 vss 0.03576f
C389 phi_fire.n5 vss 0.19603f
C390 phi_fire.t4 vss 0.0516f
C391 phi_fire.t2 vss 0.02985f
C392 phi_fire.n6 vss 0.17293f
C393 phi_fire.t8 vss 0.03833f
C394 phi_fire.n7 vss 0.11805f
C395 phi_fire.t6 vss 0.03852f
C396 phi_fire.t11 vss 0.02985f
C397 phi_fire.n8 vss 0.0392f
C398 phi_fire.t13 vss 0.03576f
C399 phi_fire.n9 vss 0.26329f
C400 phi_fire.n10 vss 0.26315f
C401 phi_fire.t3 vss 0.05223f
C402 phi_fire.n11 vss 0.40483f
C403 phi_fire.n12 vss 1.05004f
C404 phi_fire.n13 vss 0.78017f
C405 phi_fire.t1 vss 0.06015f
C406 phi_fire.n14 vss 0.25275f
C407 phi_fire.t0 vss 0.0615f
C408 vmem.t10 vss 0.07064f
C409 vmem.t9 vss 1.12982f
C410 vmem.t6 vss 0.0236f
C411 vmem.t3 vss 0.02459f
C412 vmem.n0 vss 0.02908f
C413 vmem.t11 vss 0.0152f
C414 vmem.t4 vss 0.02473f
C415 vmem.t2 vss 0.0236f
C416 vmem.n1 vss 0.04635f
C417 vmem.n2 vss 0.14042f
C418 vmem.n3 vss 0.1148f
C419 vmem.t1 vss 0.02351f
C420 vmem.t7 vss 0.02448f
C421 vmem.n4 vss 0.03065f
C422 vmem.t8 vss 0.02436f
C423 vmem.t5 vss 0.02351f
C424 vmem.n5 vss 0.02879f
C425 vmem.n6 vss 0.17627f
C426 vmem.n7 vss 0.23696f
C427 vmem.n8 vss 0.10785f
C428 vmem.t0 vss 0.01987f
C429 vdd.n0 vss 0.00406f
C430 vdd.n1 vss 0.01866f
C431 vdd.n2 vss 0.01015f
C432 vdd.n3 vss 0.00179f
C433 vdd.n4 vss 0.0078f
C434 vdd.n5 vss 0.00809f
C435 vdd.n6 vss 0.00664f
C436 vdd.n7 vss 0.0067f
C437 vdd.t43 vss 0.00251f
C438 vdd.n8 vss 0.00799f
C439 vdd.n9 vss 0.02121f
C440 vdd.n10 vss 0.00368f
C441 vdd.n11 vss 0.00248f
C442 vdd.n12 vss 0.01026f
C443 vdd.n13 vss 0.00663f
C444 vdd.n14 vss 0.00696f
C445 vdd.n15 vss 0.00431f
C446 vdd.n16 vss 0.00528f
C447 vdd.t42 vss 0.00251f
C448 vdd.n17 vss 0.00731f
C449 vdd.n18 vss 0.00231f
C450 vdd.n19 vss 0.00924f
C451 vdd.n20 vss 0.00967f
C452 vdd.n21 vss 0.0036f
C453 vdd.n22 vss 0.00602f
C454 vdd.n23 vss 0.00533f
C455 vdd.n24 vss 0.00368f
C456 vdd.n25 vss 0.01266f
C457 vdd.n26 vss 0.01143f
C458 vdd.t36 vss 0.0394f
C459 vdd.t37 vss 0
C460 vdd.n27 vss 0.02473f
C461 vdd.n28 vss 0.03939f
C462 vdd.n29 vss 0.02641f
C463 vdd.t0 vss 0.04784f
C464 vdd.n30 vss 0.03179f
C465 vdd.t9 vss 0.00307f
C466 vdd.n31 vss 0.00234f
C467 vdd.t28 vss 0.00307f
C468 vdd.t8 vss 0.02267f
C469 vdd.t44 vss 0.02267f
C470 vdd.n32 vss 0.03374f
C471 vdd.t27 vss 0.02578f
C472 vdd.n33 vss 0.03314f
C473 vdd.n34 vss 0.01819f
C474 vdd.n35 vss 0.00708f
C475 vdd.n36 vss 0.12869f
C476 vdd.t61 vss 0.00307f
C477 vdd.n37 vss 0.00234f
C478 vdd.t59 vss 0.00307f
C479 vdd.n38 vss 0.00258f
C480 vdd.t13 vss 0.00312f
C481 vdd.t58 vss 0.03959f
C482 vdd.n39 vss 0.0225f
C483 vdd.n40 vss 0.02042f
C484 vdd.t60 vss 0.04106f
C485 vdd.t47 vss 0.03405f
C486 vdd.t50 vss 0.01916f
C487 vdd.t12 vss 0.02267f
C488 vdd.n41 vss 0.01982f
C489 vdd.n42 vss 0.02923f
C490 vdd.t49 vss 0.00307f
C491 vdd.n43 vss 0.00234f
C492 vdd.t57 vss 0.00307f
C493 vdd.n44 vss 0.00258f
C494 vdd.n45 vss 0.03942f
C495 vdd.t56 vss 0.02267f
C496 vdd.t48 vss 0.02267f
C497 vdd.n46 vss 0.0318f
C498 vdd.t51 vss 0.04149f
C499 vdd.n47 vss 0.02059f
C500 vdd.t67 vss 0.00307f
C501 vdd.n48 vss 0.00258f
C502 vdd.t15 vss 0.00307f
C503 vdd.n49 vss 0.00234f
C504 vdd.t55 vss 0.00312f
C505 vdd.t17 vss 0.00312f
C506 vdd.t66 vss 0.02284f
C507 vdd.n50 vss 0.02906f
C508 vdd.n51 vss 0.02906f
C509 vdd.t14 vss 0.03242f
C510 vdd.t54 vss 0.02892f
C511 vdd.t16 vss 0.0243f
C512 vdd.t5 vss 0.02207f
C513 vdd.n52 vss 0.02041f
C514 vdd.n53 vss 0.03496f
C515 vdd.t19 vss 0.00307f
C516 vdd.n54 vss 0.00234f
C517 vdd.t24 vss 0.00307f
C518 vdd.n55 vss 0.00258f
C519 vdd.t53 vss 0.00315f
C520 vdd.t69 vss 0.00302f
C521 vdd.n56 vss 0.004f
C522 vdd.n57 vss 0.03368f
C523 vdd.t23 vss 0.02267f
C524 vdd.t18 vss 0.02267f
C525 vdd.n58 vss 0.0318f
C526 vdd.t68 vss 0.04166f
C527 vdd.t1 vss 0.02267f
C528 vdd.n59 vss 0.02041f
C529 vdd.t2 vss 0.00307f
C530 vdd.n60 vss 0.00258f
C531 vdd.t22 vss 0.00312f
C532 vdd.n61 vss 0.02162f
C533 vdd.t52 vss 0.03448f
C534 vdd.n62 vss 0.027f
C535 vdd.t4 vss 0.00312f
C536 vdd.t21 vss 0.02546f
C537 vdd.t3 vss 0.02115f
C538 vdd.n63 vss 0.03928f
C539 vdd.n64 vss 0.0043f
C540 vdd.n65 vss 0.00907f
C541 vdd.n66 vss 0.00609f
C542 vdd.n67 vss 0.00387f
C543 vdd.n68 vss 0.00747f
C544 vdd.n69 vss 0.0072f
C545 vdd.n70 vss 0.00624f
C546 vdd.n71 vss 0.00631f
C547 vdd.n72 vss 0.00361f
C548 vdd.n73 vss 0.00811f
C549 vdd.n74 vss 0.00987f
C550 vdd.n75 vss 0.00264f
C551 vdd.n76 vss 0.00565f
C552 vdd.n77 vss 0.00505f
C553 vdd.n78 vss 0.00707f
C554 vdd.n79 vss 0.00548f
C555 vdd.n80 vss 0.00279f
C556 vdd.n81 vss 0.00739f
C557 vdd.n82 vss 0.00725f
C558 vdd.n83 vss 0.00438f
C559 vdd.n84 vss 0.08015f
C560 vdd.n85 vss 0.00406f
C561 vdd.n86 vss 0.01866f
C562 vdd.n87 vss 0.00533f
C563 vdd.n88 vss 0.00179f
C564 vdd.n89 vss 0.0036f
C565 vdd.n90 vss 0.00234f
C566 vdd.n91 vss 0.00602f
C567 vdd.n92 vss 0.0132f
C568 vdd.n93 vss 0.01026f
C569 vdd.n94 vss 0.00248f
C570 vdd.n95 vss 0.0078f
C571 vdd.n96 vss 0.00368f
C572 vdd.n97 vss 0.01488f
C573 vdd.n98 vss 0.02455f
C574 vdd.t46 vss 0.00453f
C575 vdd.n99 vss 0.00739f
C576 vdd.t63 vss 0.00251f
C577 vdd.n100 vss 0.0056f
C578 vdd.n101 vss 0.00729f
C579 vdd.n102 vss 0.00617f
C580 vdd.t7 vss 0.00307f
C581 vdd.t64 vss 0.10919f
C582 vdd.t62 vss 0.10919f
C583 vdd.t45 vss 0.06135f
C584 vdd.t10 vss 0.02395f
C585 vdd.n103 vss 0.02101f
C586 vdd.t20 vss 0.02974f
C587 vdd.t6 vss 0.02816f
C588 vdd.n104 vss 0.0703f
C589 vdd.n105 vss 0.03133f
C590 vdd.n106 vss 0.0106f
C591 vdd.n107 vss 0.0427f
C592 vdd.n108 vss 0.00788f
C593 vdd.n109 vss 0.00809f
C594 vdd.n110 vss 0.00785f
C595 vdd.n111 vss 0.00928f
C596 vdd.n112 vss 0.00655f
C597 vdd.n113 vss 0.01891f
C598 vdd.n114 vss 0.00906f
C599 vdd.n115 vss 0.00347f
C600 vdd.n116 vss 0.00544f
C601 vdd.n117 vss 0.00675f
C602 vdd.n118 vss 0.00809f
C603 vdd.n119 vss 0.00969f
C604 vdd.n120 vss 0.01f
C605 vdd.t65 vss 0.00251f
C606 vdd.n121 vss 0.00735f
C607 vdd.n122 vss 0.00234f
C608 vdd.n123 vss 0.0067f
C609 vdd.n124 vss 0.00664f
C610 vdd.n125 vss 0.01015f
C611 vdd.n126 vss 0.00368f
C612 vdd.n127 vss 0.01266f
C613 vdd.n128 vss 0.01143f
C614 vdd.t33 vss 0
C615 vdd.t32 vss 0.0394f
C616 vdd.n129 vss 0.02473f
C617 vdd.n130 vss 0.03027f
C618 vdd.n131 vss 0.04766f
C619 vdd.n132 vss 0.00406f
C620 vdd.n133 vss 0.02327f
C621 vdd.n134 vss 0.01015f
C622 vdd.n135 vss 0.00179f
C623 vdd.n136 vss 0.0078f
C624 vdd.n137 vss 0.00809f
C625 vdd.n138 vss 0.00664f
C626 vdd.n139 vss 0.0067f
C627 vdd.t31 vss 0.00251f
C628 vdd.n140 vss 0.0048f
C629 vdd.t34 vss 0
C630 vdd.t35 vss 0
C631 vdd.n141 vss 0.00911f
C632 vdd.n142 vss 0.0189f
C633 vdd.n143 vss 0.01675f
C634 vdd.n144 vss 0.00368f
C635 vdd.n145 vss 0.00248f
C636 vdd.n146 vss 0.01026f
C637 vdd.n147 vss 0.00663f
C638 vdd.n148 vss 0.00696f
C639 vdd.n149 vss 0.00431f
C640 vdd.n150 vss 0.00528f
C641 vdd.t30 vss 0.00251f
C642 vdd.n151 vss 0.00731f
C643 vdd.n152 vss 0.00231f
C644 vdd.n153 vss 0.00924f
C645 vdd.n154 vss 0.00967f
C646 vdd.n155 vss 0.0036f
C647 vdd.n156 vss 0.00602f
C648 vdd.n157 vss 0.00533f
C649 vdd.n158 vss 0.00368f
C650 vdd.n159 vss 0.01675f
C651 vdd.n160 vss 0.01464f
C652 vdd.t40 vss 0
C653 vdd.t41 vss 0.00148f
C654 vdd.n161 vss 0.00933f
C655 vdd.n162 vss 0.00789f
C656 vdd.t38 vss 0.0394f
C657 vdd.t39 vss 0
C658 vdd.n163 vss 0.02473f
C659 vdd.n164 vss 0.03836f
C660 vdd.n165 vss 0.02557f
C661 vdd.t29 vss 0.02392f
C662 vdd.n166 vss 0.02101f
C663 vdd.t26 vss 0.00307f
C664 vdd.t11 vss 0.02836f
C665 vdd.t25 vss 0.029f
C666 vdd.n167 vss 0.03617f
C667 vdd.n168 vss 0.01451f
C668 vdd.n169 vss 0.05783f
C669 vdd.n170 vss 0.01135f
.ends

