* NGSPICE file created from DFF_2phase_1.ext - technology: gf180mcuD
.subckt DFF_2phase_1_pex Q D PHI_1 gated_control PHI_2 EN VDD VSS
X0 a_n1836_148# a_n2352_n394# a_n1984_n397# VSS.t20 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X1 a_972_28# a_628_148# VDD.t24 VDD.t23 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X2 VDD.t26 PHI_1.t0 a_n2820_n412# VDD.t25 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X3 a_n1984_148# D.t0 VDD.t28 VDD.t27 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X4 VDD.t7 PHI_2.t0 a_n356_n412# VDD.t6 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X5 a_n1592_n397# a_n2820_n412# a_n1836_148# VSS.t32 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X6 VSS.t12 PHI_2.t1 a_n356_n412# VSS.t11 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X7 a_872_n397# a_n356_n412# a_628_148# VSS.t17 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X8 a_n1632_148# a_n2352_n394# a_n1836_148# VDD.t20 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X9 gated_control.t1 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t1 VDD.t0 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X10 a_2093_n435# Q.t2 VSS.t14 VSS.t13 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X11 VDD.t22 a_628_148# Q.t1 VDD.t21 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X12 a_n2352_n394# a_n2820_n412# VDD.t33 VDD.t32 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X13 a_n1836_148# a_n2820_n412# a_n1984_148# VDD.t31 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X14 a_112_n394# a_n356_n412# VDD.t17 VDD.t16 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X15 a_628_148# a_n356_n412# a_480_148# VDD.t15 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X16 a_n1984_n397# D.t1 VSS.t29 VSS.t28 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X17 a_480_n397# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t9 VSS.t8 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X18 a_832_148# a_112_n394# a_628_148# VDD.t14 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X19 VDD.t30 EN.t0 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VDD.t29 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X20 a_972_28# a_628_148# VSS.t24 VSS.t23 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X21 a_n1492_28# a_n1836_148# VSS.t5 VSS.t4 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X22 gated_control.t0 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS.t1 VSS.t0 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X23 VSS.t19 a_972_28# a_872_n397# VSS.t18 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X24 a_112_n394# a_n356_n412# VSS.t16 VSS.t15 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X25 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN EN.t1 a_2093_n435# VSS.t27 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X26 VDD.t5 a_n1836_148# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t4 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X27 VSS.t7 a_n1492_28# a_n1592_n397# VSS.t6 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X28 VSS.t22 a_628_148# Q.t0 VSS.t21 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X29 VDD.t19 a_972_28# a_832_148# VDD.t18 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X30 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN Q.t3 VDD.t9 VDD.t8 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X31 VDD.t11 a_n1492_28# a_n1632_148# VDD.t10 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X32 VSS.t3 a_n1836_148# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS.t2 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X33 VSS.t26 PHI_1.t1 a_n2820_n412# VSS.t25 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X34 a_480_148# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VDD.t13 VDD.t12 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X35 a_n2352_n394# a_n2820_n412# VSS.t31 VSS.t30 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X36 a_n1492_28# a_n1836_148# VDD.t3 VDD.t2 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X37 a_628_148# a_112_n394# a_480_n397# VSS.t10 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
R0 VSS.n5 VSS.t0 2230.39
R1 VSS.t21 VSS.t23 2202.58
R2 VSS.t8 VSS.t15 2202.58
R3 VSS.t2 VSS.t4 2202.58
R4 VSS.t28 VSS.t30 2202.58
R5 VSS.n2 VSS.t2 1747.7
R6 VSS.t18 VSS.t17 1556.17
R7 VSS.t15 VSS.t11 1556.17
R8 VSS.t6 VSS.t32 1556.17
R9 VSS.t30 VSS.t25 1556.17
R10 VSS VSS.t27 1550.18
R11 VSS VSS.t21 1508.29
R12 VSS.t23 VSS.t18 1340.7
R13 VSS.t17 VSS.t10 1340.7
R14 VSS.t4 VSS.t6 1340.7
R15 VSS.t32 VSS.t20 1340.7
R16 VSS.n16 VSS 1104.92
R17 VSS.t27 VSS.t13 1101.29
R18 VSS VSS.n2 1101.29
R19 VSS.t10 VSS.t8 1005.52
R20 VSS.t20 VSS.t28 1005.52
R21 VSS.t13 VSS 700.277
R22 VSS.t0 VSS 694.292
R23 VSS.t11 VSS 694.292
R24 VSS.t25 VSS 694.292
R25 VSS.n9 VSS.t9 8.79702
R26 VSS.n14 VSS.t29 8.79702
R27 VSS.n10 VSS.n3 6.40811
R28 VSS.n15 VSS.n0 6.40811
R29 VSS.n8 VSS.n4 6.4042
R30 VSS.n13 VSS.n1 6.4042
R31 VSS.n5 VSS.t1 4.63989
R32 VSS.n7 VSS.t22 4.63989
R33 VSS.n12 VSS.t3 4.63989
R34 VSS.n6 VSS.t14 4.51271
R35 VSS.n3 VSS.t16 3.9605
R36 VSS.n0 VSS.t31 3.9605
R37 VSS.n11 VSS.n2 3.6294
R38 VSS.n4 VSS.t24 2.07392
R39 VSS.n4 VSS.t19 2.07392
R40 VSS.n1 VSS.t5 2.07392
R41 VSS.n1 VSS.t7 2.07392
R42 VSS.n3 VSS.t12 1.84987
R43 VSS.n0 VSS.t26 1.84987
R44 VSS.n9 VSS.n8 0.4385
R45 VSS.n14 VSS.n13 0.4385
R46 VSS.n8 VSS.n7 0.2965
R47 VSS.n13 VSS.n12 0.2965
R48 VSS.n6 VSS.n5 0.28
R49 VSS.n11 VSS.n10 0.2085
R50 VSS.n10 VSS.n9 0.2025
R51 VSS.n15 VSS.n14 0.2025
R52 VSS.n16 VSS 0.1645
R53 VSS.n12 VSS.n11 0.0885
R54 VSS.n7 VSS.n6 0.073
R55 VSS VSS.n16 0.047
R56 VSS VSS.n15 0.0445
R57 VDD.t21 VDD.t23 667.707
R58 VDD.t4 VDD.t2 667.707
R59 VDD.t12 VDD.t16 574.104
R60 VDD.t27 VDD.t32 574.104
R61 VDD.n5 VDD.t0 569.532
R62 VDD.n2 VDD.t4 471.139
R63 VDD VDD.t21 410.296
R64 VDD.t16 VDD.t6 405.616
R65 VDD.t32 VDD.t25 405.616
R66 VDD VDD.t29 390.017
R67 VDD.t18 VDD.t14 374.416
R68 VDD.t10 VDD.t20 374.416
R69 VDD.t29 VDD.t8 318.253
R70 VDD.t23 VDD.t18 318.253
R71 VDD.t14 VDD.t15 318.253
R72 VDD.t2 VDD.t10 318.253
R73 VDD.t20 VDD.t31 318.253
R74 VDD.n17 VDD 293.171
R75 VDD VDD.n2 288.613
R76 VDD.t15 VDD.t12 230.889
R77 VDD.t31 VDD.t27 230.889
R78 VDD.t0 VDD 195.008
R79 VDD.t6 VDD 195.008
R80 VDD.t25 VDD 195.008
R81 VDD.t8 VDD 165.368
R82 VDD.n6 VDD.t30 15.5636
R83 VDD.n15 VDD.t28 4.77854
R84 VDD.n10 VDD.t13 4.77854
R85 VDD.n12 VDD.n2 4.55932
R86 VDD.n13 VDD.t5 3.95308
R87 VDD.n8 VDD.t22 3.95308
R88 VDD.n7 VDD.t9 3.90058
R89 VDD.n5 VDD.t1 3.84351
R90 VDD.n0 VDD.t33 3.7805
R91 VDD.n3 VDD.t17 3.7805
R92 VDD.n16 VDD.n0 2.95854
R93 VDD.n14 VDD.n1 2.95854
R94 VDD.n11 VDD.n3 2.95854
R95 VDD.n9 VDD.n4 2.95854
R96 VDD.n0 VDD.t26 1.53332
R97 VDD.n3 VDD.t7 1.53332
R98 VDD.n1 VDD.t3 1.31934
R99 VDD.n1 VDD.t11 1.31934
R100 VDD.n4 VDD.t24 1.31934
R101 VDD.n4 VDD.t19 1.31934
R102 VDD.n10 VDD.n9 0.3985
R103 VDD.n15 VDD.n14 0.3985
R104 VDD.n9 VDD.n8 0.3165
R105 VDD.n14 VDD.n13 0.3165
R106 VDD.n11 VDD.n10 0.2125
R107 VDD.n16 VDD.n15 0.2125
R108 VDD.n12 VDD.n11 0.2085
R109 VDD.n7 VDD.n6 0.2045
R110 VDD.n17 VDD 0.1415
R111 VDD.n13 VDD.n12 0.0985
R112 VDD.n6 VDD.n5 0.086
R113 VDD.n8 VDD.n7 0.083
R114 VDD VDD.n16 0.0675
R115 VDD VDD.n17 0.033
R116 PHI_1.n0 PHI_1.t0 26.4265
R117 PHI_1.n0 PHI_1.t1 11.7657
R118 PHI_1 PHI_1.n0 8.04713
R119 D.n0 D.t0 29.4195
R120 D.n0 D.t1 11.4372
R121 D.n1 D 9.95
R122 D.n1 D.n0 8.0005
R123 D D.n1 0.102506
R124 PHI_2.n0 PHI_2.t0 26.4265
R125 PHI_2.n0 PHI_2.t1 11.7657
R126 PHI_2 PHI_2.n0 8.04257
R127 gated_control.n0 gated_control 16.6651
R128 gated_control.n0 gated_control.t0 4.57685
R129 gated_control gated_control.t1 4.33791
R130 gated_control gated_control.n0 0.0122931
R131 Q.n0 Q.t2 21.1948
R132 Q.n0 Q.t3 16.0605
R133 Q.n2 Q 9.45184
R134 Q Q.n1 9.13775
R135 Q.n1 Q.n0 8.12012
R136 Q.n2 Q.t0 4.5901
R137 Q Q.t1 3.91488
R138 Q Q.n2 0.150731
R139 Q.n1 Q 0.00840541
R140 EN.n0 EN.t1 19.9538
R141 EN.n0 EN.t0 17.3015
R142 EN.n1 EN 10.8498
R143 EN.n1 EN.n0 8.0005
R144 EN EN.n1 0.00742308
C0 a_628_148# VDD 0.55136f
C1 a_112_n394# PHI_1 0.01277f
C2 PHI_2 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.03773f
C3 VDD gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.34237f
C4 a_628_148# Q 0.11433f
C5 D a_n2352_n394# 0.36155f
C6 Q gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01102f
C7 a_n2820_n412# PHI_1 0.70141f
C8 EN a_n356_n412# 0.08694f
C9 PHI_2 a_2093_n435# 0
C10 a_n1836_148# a_n356_n412# 0.00268f
C11 a_112_n394# a_628_148# 0.30053f
C12 a_112_n394# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.36162f
C13 PHI_2 D 0.34149f
C14 VDD a_480_148# 0.00491f
C15 a_2093_n435# gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.0097f
C16 EN a_972_28# 0.0522f
C17 a_628_148# PHI_1 0.01804f
C18 EN a_n1492_28# 0.05124f
C19 EN gated_control 0.4397f
C20 a_n1836_148# a_n1492_28# 0.57845f
C21 a_n1836_148# gated_control 0.01329f
C22 a_n2820_n412# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00116f
C23 PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01369f
C24 PHI_2 a_480_n397# 0
C25 a_112_n394# a_480_148# 0.00294f
C26 a_n1632_148# EN 0.00368f
C27 a_872_n397# a_972_28# 0
C28 a_872_n397# gated_control 0
C29 a_n2352_n394# a_n356_n412# 0
C30 a_n1632_148# a_n1836_148# 0.01151f
C31 a_628_148# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01536f
C32 EN a_832_148# 0.00368f
C33 a_480_148# PHI_1 0.00164f
C34 VDD EN 0.35601f
C35 PHI_2 a_n356_n412# 0.60119f
C36 VDD a_n1836_148# 0.56047f
C37 a_n1492_28# a_n2352_n394# 0.00888f
C38 a_n2352_n394# gated_control 0.00668f
C39 EN Q 0.38669f
C40 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_n356_n412# 0
C41 a_628_148# a_480_148# 0
C42 a_n1984_n397# EN 0.0022f
C43 a_112_n394# EN 0.05124f
C44 a_n1984_n397# a_n1836_148# 0
C45 PHI_2 a_972_28# 0.03174f
C46 PHI_2 a_n1492_28# 0.03207f
C47 PHI_2 gated_control 0.31085f
C48 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN gated_control 0.33472f
C49 a_n2820_n412# EN 0.08666f
C50 EN PHI_1 0.059f
C51 a_n2820_n412# a_n1836_148# 0.07055f
C52 a_n1836_148# PHI_1 0.01882f
C53 PHI_2 a_n1632_148# 0.00411f
C54 VDD a_n2352_n394# 0.4225f
C55 VDD a_n1984_148# 0.00491f
C56 PHI_2 a_832_148# 0.00422f
C57 a_2093_n435# gated_control 0.00113f
C58 a_n1592_n397# EN 0.00577f
C59 PHI_2 VDD 0.46604f
C60 a_628_148# EN 0.11443f
C61 a_n1592_n397# a_n1836_148# 0.01595f
C62 D a_n1492_28# 0.00242f
C63 a_n1984_n397# a_n2352_n394# 0.00194f
C64 D gated_control 0.17162f
C65 EN gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.20415f
C66 PHI_2 Q 0.32019f
C67 a_n1836_148# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.09501f
C68 VDD gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.42344f
C69 PHI_2 a_n1984_n397# 0
C70 a_628_148# a_872_n397# 0.01595f
C71 a_n2820_n412# a_n2352_n394# 0.30528f
C72 PHI_2 a_112_n394# 0.07395f
C73 Q gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08537f
C74 a_n2352_n394# PHI_1 0.0533f
C75 gated_control a_480_n397# 0
C76 EN a_480_148# 0.00101f
C77 a_n1984_148# PHI_1 0.00201f
C78 a_112_n394# gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C79 PHI_2 a_n2820_n412# 0.02723f
C80 D VDD 0.18262f
C81 Q a_2093_n435# 0.00241f
C82 PHI_2 PHI_1 2.45879f
C83 a_972_28# a_n356_n412# 0.02403f
C84 a_n2352_n394# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C85 a_n1492_28# a_n356_n412# 0
C86 gated_control a_n356_n412# 0.00985f
C87 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.01636f
C88 PHI_2 a_n1592_n397# 0
C89 a_n1984_n397# D 0
C90 PHI_2 a_628_148# 0.04011f
C91 PHI_2 gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.45413f
C92 a_628_148# gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C93 a_972_28# gated_control 0.01014f
C94 a_n1492_28# gated_control 0.00972f
C95 D a_n2820_n412# 0.15891f
C96 D PHI_1 0.0221f
C97 a_n1836_148# EN 0.11055f
C98 a_112_n394# a_480_n397# 0.00194f
C99 VDD a_n356_n412# 1.03607f
C100 PHI_2 a_480_148# 0
C101 a_n1632_148# a_n1492_28# 0.00109f
C102 a_n1632_148# gated_control 0
C103 a_872_n397# EN 0.00579f
C104 Q a_n356_n412# 0.00225f
C105 a_972_28# a_832_148# 0.00109f
C106 gated_control a_832_148# 0
C107 D gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.01068f
C108 VDD a_972_28# 0.32599f
C109 a_112_n394# a_n356_n412# 0.30528f
C110 VDD a_n1492_28# 0.32599f
C111 VDD gated_control 0.26726f
C112 Q a_972_28# 0.25874f
C113 EN a_n2352_n394# 0.05107f
C114 Q gated_control 0.22358f
C115 a_628_148# a_480_n397# 0
C116 a_n1836_148# a_n2352_n394# 0.30053f
C117 a_n2820_n412# a_n356_n412# 0
C118 a_480_n397# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0
C119 PHI_1 a_n356_n412# 0.01733f
C120 VDD a_n1632_148# 0.01506f
C121 EN a_n1984_148# 0.00101f
C122 a_n1836_148# a_n1984_148# 0
C123 a_n1984_n397# gated_control 0
C124 a_112_n394# a_972_28# 0.00888f
C125 a_112_n394# gated_control 0.00668f
C126 PHI_2 EN 0.1362f
C127 VDD a_832_148# 0.01506f
C128 PHI_2 a_n1836_148# 0.04895f
C129 a_n2820_n412# a_n1492_28# 0.02403f
C130 a_972_28# PHI_1 0.01261f
C131 a_628_148# a_n356_n412# 0.07055f
C132 a_n2820_n412# gated_control 0.00985f
C133 EN gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.65271f
C134 a_n1492_28# PHI_1 0.01314f
C135 gated_control PHI_1 0.00846f
C136 gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q a_n356_n412# 0.16689f
C137 VDD Q 0.37581f
C138 PHI_2 a_872_n397# 0
C139 EN a_2093_n435# 0.00398f
C140 a_112_n394# VDD 0.42245f
C141 a_n1632_148# PHI_1 0.00534f
C142 a_n1592_n397# a_n1492_28# 0
C143 a_628_148# a_972_28# 0.57845f
C144 a_n1592_n397# gated_control 0
C145 a_n2352_n394# a_n1984_148# 0.00294f
C146 a_628_148# gated_control 0.01553f
C147 D EN 0.13355f
C148 a_972_28# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.00242f
C149 a_n1492_28# gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.2556f
C150 a_112_n394# Q 0.00101f
C151 gated_control gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q 0.23535f
C152 PHI_1 a_832_148# 0.00477f
C153 D a_n1836_148# 0.01538f
C154 PHI_2 a_n2352_n394# 0.03321f
C155 VDD a_n2820_n412# 0.99732f
C156 VDD PHI_1 0.98251f
C157 PHI_2 a_n1984_148# 0
C158 Q PHI_1 0.03331f
C159 EN a_480_n397# 0.0022f
C160 a_628_148# a_832_148# 0.01151f
C161 gated_control VSS 1.67727f
C162 EN VSS 2.71676f
C163 Q VSS 1.01402f
C164 PHI_2 VSS 2.77872f
C165 D VSS 0.48547f
C166 PHI_1 VSS 3.51163f
C167 VDD VSS 13.6464f
C168 a_2093_n435# VSS 0.0072f
C169 a_480_n397# VSS 0.0042f
C170 a_872_n397# VSS 0.0095f
C171 gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN VSS 0.77496f
C172 a_n1984_n397# VSS 0.0042f
C173 a_n1592_n397# VSS 0.0095f
C174 a_972_28# VSS 0.42076f
C175 a_112_n394# VSS 0.53018f
C176 a_628_148# VSS 1.13543f
C177 gf180mcu_fd_sc_mcu9t5v0__latq_1_1.Q VSS 0.66898f
C178 a_n1492_28# VSS 0.42076f
C179 a_n2352_n394# VSS 0.53018f
C180 a_n356_n412# VSS 1.18728f
C181 a_n1836_148# VSS 1.14251f
C182 a_n2820_n412# VSS 1.19329f
C183 PHI_2.t0 VSS 0.09365f
C184 PHI_2.t1 VSS 0.05178f
C185 PHI_2.n0 VSS 0.09322f
C186 PHI_1.t0 VSS 0.09191f
C187 PHI_1.t1 VSS 0.05082f
C188 PHI_1.n0 VSS 0.09144f
.ends

