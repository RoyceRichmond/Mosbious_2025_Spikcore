* Extracted by KLayout with GF180MCU LVS runset on : 28/07/2025 08:10

.SUBCKT DFF_2phase_1 VSS|vss D|Q|out_m Q|q E|phi_2 VDD|vdd D E|phi_1 vss
M$1 VDD|vdd E|phi_2 \$2 \$21 pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$2 \$3 \$2 VDD|vdd \$21 pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$3 \$24 D|Q|out_m VDD|vdd \$21 pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$4 \$5 \$2 \$24 \$21 pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U PD=1.52U
M$5 \$5 \$3 \$23 \$21 pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U PD=1.52U
M$6 VDD|vdd \$6 \$23 \$21 pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$7 \$6 \$5 VDD|vdd \$21 pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$8 VDD|vdd \$5 Q|q \$21 pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$9 VDD|vdd E|phi_1 \$17 \$41 pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$10 \$18 \$17 VDD|vdd \$41 pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$11 \$36 D VDD|vdd \$41 pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$12 \$27 \$17 \$36 \$41 pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$13 \$27 \$18 \$37 \$41 pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$14 VDD|vdd \$28 \$37 \$41 pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$15 \$28 \$27 VDD|vdd \$41 pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$16 VDD|vdd \$27 D|Q|out_m \$41 pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$17 \$9 D|Q|out_m VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$18 \$5 \$3 \$9 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$19 \$11 \$2 \$5 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$20 VSS|vss \$6 \$11 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$21 \$6 \$5 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$22 VSS|vss E|phi_2 \$2 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$23 \$3 \$2 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$24 VSS|vss \$5 Q|q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$25 \$30 D VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$26 \$27 \$18 \$30 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$27 \$34 \$17 \$27 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$28 VSS|vss \$28 \$34 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$29 \$28 \$27 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$30 VSS|vss E|phi_1 \$17 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$31 \$18 \$17 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$32 VSS|vss \$27 D|Q|out_m vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
.ENDS DFF_2phase_1
