magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l33d0 >>
<< l34d0 >>
<< l30d0 >>
<< l22d0 >>
<< l31d0 >>
<< l32d0 >>
<< labels >>
rlabel l34d10 -0.092 0.0065 -0.092 0.0065 0 
<< end >>
