* NGSPICE file created from swmatrix_row_10.ext - technology: gf180mcuD

.subckt swmatrix_row_10_pex D_out D_in PHI_1 PHI_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] VDD
+ pin VSS
X0 pin.t52 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 BUS[7].t16 vdd.t85 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X1 pin.t187 swmatrix_Tgate_8.gated_control BUS[2].t21 vss.t301 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X2 swmatrix_Tgate_3.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t91 vdd.t90 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 BUS[7].t15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t51 vdd.t84 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X4 BUS[1].t17 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 pin.t197 vdd.t401 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X5 vdd.t518 a_51256_2002# a_51116_2122# vdd.t517 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X6 a_26296_2002# a_25952_2122# vss.t360 vss.t359 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X7 BUS[5].t23 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 pin.t154 vdd.t332 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X8 a_34508_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t259 vss.t258 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X9 a_53620_1577# a_52392_1562# a_53376_2122# vss.t190 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X10 a_6716_1580# a_6248_1562# vss.t45 vss.t44 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X11 BUS[6].t23 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 pin.t102 vdd.t237 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X12 BUS[4].t17 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 pin.t60 vdd.t154 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X13 vdd.t224 PHI_2.t0 a_39912_1562# vdd.t223 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X14 BUS[8].t10 swmatrix_Tgate_3.gated_control pin.t107 vss.t214 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X15 a_4921_1539# ShiftReg_row_10_2$1_0.Q[1] vss.t81 vss.t80 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X16 pin.t19 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 BUS[8].t4 vdd.t43 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X17 vdd.t22 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t21 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X18 pin.t121 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 BUS[6].t22 vdd.t258 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X19 BUS[9].t14 swmatrix_Tgate_1.gated_control pin.t196 vss.t311 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X20 pin.t79 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 BUS[4].t16 vdd.t212 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X21 vss.t283 a_45016_2002# a_44916_1577# vss.t282 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X22 vdd.t186 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] vdd.t185 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X23 vss.t321 a_38776_2002# a_38676_1577# vss.t320 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X24 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t0 a_11161_1539# vss.t184 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X25 a_44156_1580# a_43688_1562# vss.t187 vss.t186 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X26 a_13472_2122# a_12488_1562# a_13324_2122# vdd.t67 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X27 a_19564_2122# ShiftReg_row_10_2$1_0.Q[3] vdd.t167 vdd.t166 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X28 vdd.t263 a_53720_2002# a_53580_2122# vdd.t262 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X29 vss.t234 PHI_1.t0 a_56168_1562# vss.t233 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X30 BUS[8].t22 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t235 vdd.t531 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X31 vdd.t509 enable.t1 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t508 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X32 pin.t195 swmatrix_Tgate_1.gated_control BUS[9].t13 vss.t310 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X33 a_26156_2122# a_25436_1580# a_25952_2122# vdd.t147 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X34 a_56636_1580# a_56168_1562# vdd.t501 vdd.t500 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X35 a_19916_2122# a_19196_1580# a_19712_2122# vdd.t387 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X36 swmatrix_Tgate_7.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t37 vdd.t36 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X37 BUS[7].t14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 pin.t50 vdd.t83 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X38 vdd.t286 PHI_1.t1 a_12488_1562# vdd.t285 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X39 BUS[4].t23 swmatrix_Tgate_7.gated_control pin.t224 vss.t389 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X40 pin.t202 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 BUS[9].t16 vdd.t421 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X41 BUS[5].t5 swmatrix_Tgate_5.gated_control pin.t8 vss.t19 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X42 a_7576_2002# a_7232_2122# vdd.t443 vdd.t442 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X43 pin.t49 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[7].t23 vdd.t82 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X44 swmatrix_Tgate_2.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t503 vdd.t502 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X45 swmatrix_Tgate_1.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t244 vss.t243 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X46 vss.t377 a_47480_2002# a_47380_1577# vss.t376 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X47 vdd.t288 PHI_1.t2 a_8_1562# vdd.t287 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X48 vss.t28 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t27 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X49 pin.t80 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 BUS[4].t15 vdd.t213 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X50 BUS[2].t8 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 pin.t159 vdd.t341 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X51 a_48601_1539# ShiftReg_row_10_2$1_0.Q[8] vss.t168 vss.t167 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X52 a_46620_1580# a_46152_1562# vss.t57 vss.t56 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X53 vss.t192 PHI_2.t1 a_58632_1562# vss.t191 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X54 a_34900_1577# a_33672_1562# a_34656_2122# vss.t257 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X55 pin.t7 swmatrix_Tgate_5.gated_control BUS[5].t4 vss.t18 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X56 a_28620_2122# a_27900_1580# a_28416_2122# vdd.t168 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X57 BUS[6].t21 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 pin.t122 vdd.t259 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X58 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[5] vdd.t133 vdd.t132 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X59 vss.t254 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t253 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X60 vss.t358 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t357 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X61 a_45016_2002# a_44672_2122# vdd.t16 vdd.t15 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X62 vss.t242 PHI_1.t3 a_8_1562# vss.t241 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X63 BUS[7].t5 swmatrix_Tgate_0.gated_control pin.t25 vss.t54 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X64 pin.t123 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[6].t20 vdd.t260 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X65 vdd.t108 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t107 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X66 vss.t194 PHI_2.t2 a_2472_1562# vss.t193 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X67 vdd.t412 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t411 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X68 pin.t127 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 BUS[3].t17 vdd.t278 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X69 a_32044_2122# ShiftReg_row_10_2$1_0.Q[5] vdd.t131 vdd.t130 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X70 vss.t300 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t299 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X71 vss.t204 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t203 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X72 a_2940_1580# a_2472_1562# vdd.t113 vdd.t112 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X73 pin.t48 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 BUS[7].t22 vdd.t81 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X74 pin.t228 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 BUS[10].t23 vdd.t498 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X75 a_53376_2122# a_52860_1580# a_53228_1577# vss.t249 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X76 pin.t219 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 BUS[2].t22 vdd.t487 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X77 vdd.t104 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t103 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X78 swmatrix_Tgate_5.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t7 vss.t6 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X79 BUS[9].t17 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t203 vdd.t422 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X80 a_28760_2002# a_28416_2122# vss.t330 vss.t329 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X81 BUS[7].t21 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t47 vdd.t80 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X82 BUS[1].t16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t198 vdd.t402 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X83 a_47480_2002# a_47136_2122# vdd.t124 vdd.t123 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X84 vss.t143 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] vss.t142 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X85 BUS[5].t22 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t100 vdd.t235 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X86 a_23641_1539# ShiftReg_row_10_2$1_0.Q[4] vss.t315 vss.t314 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X87 vss.t196 PHI_2.t3 a_39912_1562# vss.t195 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X88 a_7084_1577# ShiftReg_row_10_2$1_0.Q[1] vss.t79 vss.t78 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X89 a_1336_2002# a_992_2122# vss.t115 vss.t114 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X90 vdd.t462 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] vdd.t461 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X91 pin.t176 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 BUS[9].t7 vdd.t358 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X92 BUS[3].t23 swmatrix_Tgate_4.gated_control pin.t53 vss.t106 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X93 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[2] vdd.t447 vdd.t446 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X94 vdd.t437 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] vdd.t436 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X95 pin.t111 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 BUS[1].t15 vdd.t244 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X96 a_61081_1539# d_out.t2 vss.t335 vss.t334 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X97 pin.t221 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 BUS[3].t16 vdd.t491 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X98 a_27900_1580# a_27432_1562# vss.t375 vss.t374 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X99 vss.t309 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t308 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X100 pin.t12 swmatrix_Tgate_5.gated_control BUS[5].t3 vss.t17 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X101 vdd.t138 a_59616_2122# d_out.t1 vdd.t137 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X102 a_32192_2122# a_31676_1580# a_32044_1577# vss.t92 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X103 a_25952_2122# a_25436_1580# a_25804_1577# vss.t144 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X104 BUS[3].t15 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 pin.t63 vdd.t187 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X105 a_44524_1577# ShiftReg_row_10_2$1_0.Q[7] vss.t355 vss.t354 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X106 pin.t30 swmatrix_Tgate_6.gated_control BUS[6].t5 vss.t74 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X107 vdd.t280 PHI_1.t4 a_49928_1562# vdd.t279 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X108 pin.t227 swmatrix_Tgate_7.gated_control BUS[4].t22 vss.t388 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X109 vdd.t511 enable.t2 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t510 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X110 BUS[8].t23 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 pin.t236 vdd.t532 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X111 vdd.t513 enable.t3 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t512 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X112 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t4 a_48601_1539# vss.t41 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X113 vss.t236 PHI_1.t5 a_12488_1562# vss.t235 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X114 BUS[2].t23 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 pin.t220 vdd.t488 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X115 a_59468_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t398 vdd.t397 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X116 a_53376_2122# a_52392_1562# a_53228_2122# vdd.t197 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X117 pin.t101 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 BUS[5].t21 vdd.t236 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X118 a_12956_1580# a_12488_1562# vdd.t66 vdd.t65 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X119 a_22520_2002# a_22176_2122# vdd.t460 vdd.t459 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X120 BUS[8].t9 swmatrix_Tgate_3.gated_control pin.t106 vss.t213 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X121 BUS[6].t4 swmatrix_Tgate_6.gated_control pin.t29 vss.t73 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X122 pin.t217 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[8].t20 vdd.t485 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X123 pin.t81 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[4].t14 vdd.t214 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X124 pin.t174 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[2].t14 vdd.t356 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X125 a_45016_2002# a_44672_2122# vss.t11 vss.t10 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X126 vss.t16 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t15 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X127 a_46988_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t30 vss.t29 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X128 pin.t105 swmatrix_Tgate_3.gated_control BUS[8].t8 vss.t212 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X129 a_41240_2002# a_40896_2122# vss.t381 vss.t380 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X130 a_844_2122# D_in.t0 vdd.t294 vdd.t293 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X131 vss.t149 a_10040_2002# a_9940_1577# vss.t148 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X132 BUS[1].t14 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 pin.t112 vdd.t245 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X133 vdd.t32 PHI_2.t4 a_52392_1562# vdd.t31 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X134 BUS[4].t13 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t114 vdd.t247 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X135 vss.t35 PHI_2.t5 a_21192_1562# vss.t34 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X136 vdd.t449 a_35000_2002# a_34860_2122# vdd.t448 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X137 swmatrix_Tgate_9.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t470 vdd.t469 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X138 a_21660_1580# a_21192_1562# vdd.t30 vdd.t29 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X139 vss.t341 a_57496_2002# a_57396_1577# vss.t340 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X140 a_38284_2122# ShiftReg_row_10_2$1_0.Q[6] vdd.t180 vdd.t179 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X141 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[1] vdd.t89 vdd.t88 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X142 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t5 a_23641_1539# vss.t42 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X143 a_32192_2122# a_31208_1562# a_32044_2122# vdd.t142 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X144 pin.t218 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 BUS[8].t21 vdd.t486 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X145 a_56636_1580# a_56168_1562# vss.t392 vss.t391 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X146 a_9180_1580# a_8712_1562# vdd.t383 vdd.t382 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X147 a_25952_2122# a_24968_1562# a_25804_2122# vdd.t516 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X148 a_34508_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t340 vdd.t339 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X149 a_44916_1577# a_43688_1562# a_44672_2122# vss.t185 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X150 a_38636_2122# a_37916_1580# a_38432_2122# vdd.t316 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X151 BUS[10].t22 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 pin.t164 vdd.t346 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X152 a_25804_1577# ShiftReg_row_10_2$1_0.Q[4] vss.t313 vss.t312 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X153 BUS[8].t2 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t5 vdd.t19 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X154 vss.t3 a_1336_2002# a_1236_1577# vss.t2 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X155 a_20056_2002# a_19712_2122# vss.t409 vss.t408 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X156 BUS[4].t12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t115 vdd.t248 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X157 a_22028_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t164 vss.t163 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X158 a_16180_1577# a_14952_1562# a_15936_2122# vss.t230 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X159 pin.t132 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 BUS[10].t21 vdd.t297 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X160 a_9548_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t147 vss.t146 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X161 pin.t85 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 BUS[6].t19 vdd.t218 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X162 pin.t116 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[4].t11 vdd.t249 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X163 pin.t177 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[9].t8 vdd.t359 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X164 vss.t105 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t104 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X165 a_47340_2122# a_46620_1580# a_47136_2122# vdd.t139 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X166 a_22520_2002# a_22176_2122# vss.t364 vss.t363 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X167 BUS[2].t15 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t175 vdd.t357 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X168 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[8] vdd.t174 vdd.t173 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X169 a_13324_2122# ShiftReg_row_10_2$1_0.Q[2] vdd.t445 vdd.t444 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X170 vss.t9 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t8 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X171 vss.t5 a_3800_2002# a_3700_1577# vss.t4 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X172 vdd.t34 PHI_2.t6 a_33672_1562# vdd.t33 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X173 pin.t24 swmatrix_Tgate_0.gated_control BUS[7].t4 vss.t53 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X174 vss.t238 PHI_1.t6 a_49928_1562# vss.t237 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X175 a_28416_2122# a_27900_1580# a_28268_1577# vss.t162 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X176 BUS[9].t0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t59 vdd.t118 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X177 a_57496_2002# a_57152_2122# vdd.t378 vdd.t377 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X178 a_2940_1580# a_2472_1562# vss.t111 vss.t110 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X179 vdd.t373 a_16280_2002# a_16140_2122# vdd.t372 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X180 vdd.t320 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t319 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X181 pin.t124 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 BUS[2].t0 vdd.t261 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X182 vdd.t458 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t457 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X183 a_50764_2122# ShiftReg_row_10_2$1_0.Q[8] vdd.t172 vdd.t171 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X184 BUS[1].t23 swmatrix_Tgate_9.gated_control pin.t99 vss.t202 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X185 a_19196_1580# a_18728_1562# vdd.t161 vdd.t160 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X186 a_7476_1577# a_6248_1562# a_7232_2122# vss.t43 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X187 BUS[3].t22 swmatrix_Tgate_4.gated_control pin.t57 vss.t103 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X188 pin.t46 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[7].t20 vdd.t79 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X189 a_37916_1580# a_37448_1562# vss.t225 vss.t224 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X190 pin.t0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[5].t20 vdd.t8 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X191 pin.t64 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 BUS[3].t14 vdd.t188 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X192 a_15788_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t371 vdd.t370 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X193 a_1336_2002# a_992_2122# vdd.t117 vdd.t116 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X194 pin.t98 swmatrix_Tgate_9.gated_control BUS[1].t22 vss.t201 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X195 swmatrix_Tgate_0.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t227 vss.t226 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X196 BUS[10].t20 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 pin.t133 vdd.t298 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X197 vss.t370 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] vss.t369 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X198 pin.t56 swmatrix_Tgate_4.gated_control BUS[3].t21 vss.t102 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X199 BUS[1].t13 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t113 vdd.t246 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X200 a_42361_1539# ShiftReg_row_10_2$1_0.Q[7] vss.t353 vss.t352 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X201 swmatrix_Tgate_4.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t97 vdd.t96 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X202 BUS[5].t19 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t1 vdd.t9 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X203 BUS[9].t20 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t214 vdd.t479 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X204 vdd.t146 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] vdd.t145 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X205 vdd.t429 a_7576_2002# a_7436_2122# vdd.t428 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X206 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[4] vdd.t407 vdd.t406 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X207 a_9940_1577# a_8712_1562# a_9696_2122# vss.t286 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X208 vdd.t39 enable.t6 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t38 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X209 vss.t345 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t344 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X210 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN d_out.t3 vdd.t431 vdd.t430 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X211 a_44672_2122# a_44156_1580# a_44524_1577# vss.t46 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X212 vss.t176 a_20056_2002# a_19956_1577# vss.t175 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X213 a_28416_2122# a_27432_1562# a_28268_2122# vdd.t483 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X214 vss.t66 a_13816_2002# a_13716_1577# vss.t65 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X215 pin.t23 swmatrix_Tgate_0.gated_control BUS[7].t3 vss.t52 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X216 a_12956_1580# a_12488_1562# vss.t77 vss.t76 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X217 vss.t240 PHI_1.t7 a_31208_1562# vss.t239 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X218 BUS[1].t12 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t143 vdd.t312 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X219 vdd.t380 a_45016_2002# a_44876_2122# vdd.t379 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X220 BUS[5].t18 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t2 vdd.t10 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X221 a_28268_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t124 vss.t123 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X222 a_38776_2002# a_38432_2122# vdd.t366 vdd.t365 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X223 BUS[3].t13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t61 vdd.t162 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X224 BUS[10].t19 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 pin.t77 vdd.t210 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X225 a_31676_1580# a_31208_1562# vdd.t141 vdd.t140 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X226 a_41240_2002# a_40896_2122# vdd.t495 vdd.t494 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X227 pin.t144 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[1].t11 vdd.t313 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X228 pin.t26 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[5].t17 vdd.t60 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X229 BUS[8].t7 swmatrix_Tgate_3.gated_control pin.t110 vss.t211 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X230 a_57496_2002# a_57152_2122# vss.t281 vss.t280 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X231 a_59960_2002# a_59616_2122# vss.t135 vss.t134 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X232 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t7 a_4921_1539# vss.t181 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X233 vss.t117 a_22520_2002# a_22420_1577# vss.t116 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X234 pin.t65 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[4].t10 vdd.t198 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X235 a_21660_1580# a_21192_1562# vss.t33 vss.t32 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X236 pin.t16 swmatrix_Tgate_2.gated_control BUS[10].t5 vss.t26 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X237 vss.t37 PHI_2.t7 a_33672_1562# vss.t36 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X238 BUS[8].t3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 pin.t6 vdd.t20 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X239 a_40380_1580# a_39912_1562# vdd.t369 vdd.t368 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X240 BUS[6].t18 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t86 vdd.t219 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X241 a_9180_1580# a_8712_1562# vss.t285 vss.t284 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X242 a_26196_1577# a_24968_1562# a_25952_2122# vss.t397 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X243 BUS[4].t9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 pin.t66 vdd.t199 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X244 a_19956_1577# a_18728_1562# a_19712_2122# vss.t157 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X245 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t8 a_42361_1539# vss.t182 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X246 a_7232_2122# a_6716_1580# a_7084_1577# vss.t356 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X247 BUS[2].t20 swmatrix_Tgate_8.gated_control pin.t186 vss.t298 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X248 a_20056_2002# a_19712_2122# vdd.t536 vdd.t535 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X249 a_53228_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t106 vdd.t105 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X250 a_44672_2122# a_43688_1562# a_44524_2122# vdd.t194 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X251 pin.t206 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[8].t11 vdd.t463 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X252 vdd.t190 enable.t9 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t189 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X253 pin.t87 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[6].t17 vdd.t220 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X254 a_57356_2122# a_56636_1580# a_57152_2122# vdd.t415 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X255 pin.t45 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[7].t19 vdd.t78 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X256 swmatrix_Tgate_1.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t290 vdd.t289 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X257 swmatrix_Tgate_3.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t83 vss.t82 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X258 pin.t185 swmatrix_Tgate_8.gated_control BUS[2].t19 vss.t297 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X259 a_3800_2002# a_3456_2122# vdd.t184 vdd.t183 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X260 BUS[10].t18 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 pin.t78 vdd.t211 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X261 BUS[1].t10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 pin.t145 vdd.t314 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X262 a_32536_2002# a_32192_2122# vss.t252 vss.t251 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X263 BUS[5].t16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 pin.t27 vdd.t61 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X264 a_40748_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t108 vss.t107 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X265 vdd.t282 PHI_1.t8 a_43688_1562# vdd.t281 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X266 vdd.t476 a_26296_2002# a_26156_2122# vdd.t475 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X267 a_9696_2122# a_9180_1580# a_9548_1577# vss.t145 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X268 BUS[9].t21 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 pin.t215 vdd.t480 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X269 a_28660_1577# a_27432_1562# a_28416_2122# vss.t373 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X270 a_59100_1580# a_58632_1562# vdd.t394 vdd.t393 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X271 a_1196_2122# a_476_1580# a_992_2122# vdd.t23 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X272 vss.t87 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] vss.t86 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X273 pin.t44 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[7].t18 vdd.t77 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X274 pin.t152 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[1].t9 vdd.t330 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X275 pin.t166 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 BUS[2].t10 vdd.t348 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X276 vdd.t255 PHI_2.t8 a_14952_1562# vdd.t254 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X277 a_476_1580# a_8_1562# vdd.t54 vdd.t53 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X278 pin.t207 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[8].t12 vdd.t464 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X279 pin.t204 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[9].t18 vdd.t432 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X280 pin.t88 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[6].t16 vdd.t221 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X281 a_59820_2122# a_59100_1580# a_59616_2122# vdd.t57 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X282 a_25804_2122# ShiftReg_row_10_2$1_0.Q[4] vdd.t405 vdd.t404 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X283 pin.t97 swmatrix_Tgate_9.gated_control BUS[1].t21 vss.t200 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X284 a_47136_2122# a_46620_1580# a_46988_1577# vss.t136 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X285 BUS[10].t17 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 pin.t200 vdd.t408 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X286 a_19196_1580# a_18728_1562# vss.t156 vss.t155 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X287 BUS[8].t13 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t208 vdd.t465 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X288 vdd.t99 a_28760_2002# a_28620_2122# vdd.t98 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X289 BUS[6].t15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 pin.t89 vdd.t222 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X290 a_7232_2122# a_6248_1562# a_7084_2122# vdd.t42 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X291 pin.t194 swmatrix_Tgate_1.gated_control BUS[9].t12 vss.t307 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X292 vdd.t14 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t13 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X293 a_3660_2122# a_2940_1580# a_3456_2122# vdd.t134 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X294 pin.t162 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 BUS[10].t16 vdd.t344 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X295 vdd.t46 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vdd.t45 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X296 BUS[4].t21 swmatrix_Tgate_7.gated_control pin.t226 vss.t387 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X297 vss.t113 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t112 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X298 vss.t126 a_59960_2002# a_59860_1577# vss.t125 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X299 vdd.t284 PHI_1.t9 a_6248_1562# vdd.t283 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X300 swmatrix_Tgate_2.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t394 vss.t393 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X301 pin.t205 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[9].t19 vdd.t433 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X302 pin.t43 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 BUS[7].t17 vdd.t76 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X303 swmatrix_Tgate_6.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t51 vdd.t50 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X304 a_54841_1539# ShiftReg_row_10_2$1_0.Q[9] vss.t326 vss.t325 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X305 a_9696_2122# a_8712_1562# a_9548_2122# vdd.t381 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X306 BUS[2].t11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 pin.t167 vdd.t349 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X307 a_41100_2122# a_40380_1580# a_40896_2122# vdd.t35 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X308 pin.t11 swmatrix_Tgate_5.gated_control BUS[5].t2 vss.t14 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X309 BUS[9].t4 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t160 vdd.t342 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X310 vdd.t474 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] vdd.t473 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X311 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[7] vdd.t453 vdd.t452 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X312 BUS[7].t12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t42 vdd.t75 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X313 a_19712_2122# a_19196_1580# a_19564_1577# vss.t290 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X314 pin.t135 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[2].t2 vdd.t300 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X315 a_3800_2002# a_3456_2122# vss.t180 vss.t179 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X316 vdd.t152 a_10040_2002# a_9900_2122# vdd.t151 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X317 BUS[7].t2 swmatrix_Tgate_0.gated_control pin.t22 vss.t51 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X318 a_59100_1580# a_58632_1562# vss.t293 vss.t292 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X319 vdd.t257 PHI_2.t9 a_8712_1562# vdd.t256 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X320 a_47136_2122# a_46152_1562# a_46988_2122# vdd.t49 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X321 vss.t170 a_32536_2002# a_32436_1577# vss.t169 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X322 pin.t62 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 BUS[3].t12 vdd.t163 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X323 a_1236_1577# a_8_1562# a_992_2122# vss.t62 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X324 pin.t163 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[10].t15 vdd.t345 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X325 a_31676_1580# a_31208_1562# vss.t139 vss.t138 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X326 vdd.t441 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t440 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X327 BUS[8].t14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t209 vdd.t466 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X328 vss.t248 PHI_1.t10 a_43688_1562# vss.t247 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X329 a_38776_2002# a_38432_2122# vss.t269 vss.t268 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X330 BUS[5].t15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 pin.t28 vdd.t62 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X331 a_59960_2002# a_59616_2122# vdd.t136 vdd.t135 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X332 a_50396_1580# a_49928_1562# vdd.t386 vdd.t385 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X333 pin.t109 swmatrix_Tgate_3.gated_control BUS[8].t6 vss.t210 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X334 BUS[3].t11 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 pin.t199 vdd.t403 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X335 a_53720_2002# a_53376_2122# vdd.t472 vdd.t471 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X336 a_13676_2122# a_12956_1580# a_13472_2122# vdd.t191 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X337 BUS[9].t5 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t168 vdd.t350 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X338 BUS[10].t14 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t130 vdd.t295 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X339 BUS[7].t11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 pin.t41 vdd.t74 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X340 swmatrix_Tgate_8.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t243 vdd.t242 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X341 BUS[4].t8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t67 vdd.t200 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X342 vss.t218 PHI_2.t10 a_14952_1562# vss.t217 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X343 vdd.t64 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t63 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X344 vdd.t5 a_1336_2002# a_1196_2122# vdd.t4 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X345 pin.t169 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[9].t6 vdd.t351 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X346 vss.t154 a_41240_2002# a_41140_1577# vss.t153 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X347 a_15420_1580# a_14952_1562# vdd.t271 vdd.t270 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X348 pin.t153 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 BUS[1].t8 vdd.t331 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X349 pin.t68 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 BUS[4].t7 vdd.t201 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X350 a_40380_1580# a_39912_1562# vss.t272 vss.t271 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X351 vss.t220 PHI_2.t11 a_52392_1562# vss.t219 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X352 a_19712_2122# a_18728_1562# a_19564_2122# vdd.t159 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X353 a_22380_2122# a_21660_1580# a_22176_2122# vdd.t374 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X354 BUS[5].t14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t125 vdd.t276 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X355 a_52860_1580# a_52392_1562# vdd.t196 vdd.t195 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X356 a_38676_1577# a_37448_1562# a_38432_2122# vss.t223 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X357 BUS[6].t14 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t118 vdd.t251 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X358 BUS[3].t10 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 pin.t155 vdd.t333 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X359 vss.t407 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t406 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X360 pin.t225 swmatrix_Tgate_7.gated_control BUS[4].t20 vss.t386 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X361 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t10 a_61081_1539# vss.t205 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X362 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t11 a_54841_1539# vss.t206 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X363 a_19564_1577# ShiftReg_row_10_2$1_0.Q[3] vss.t161 vss.t160 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X364 vdd.t305 PHI_1.t11 a_24968_1562# vdd.t304 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X365 a_32536_2002# a_32192_2122# vdd.t318 vdd.t317 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X366 BUS[2].t18 swmatrix_Tgate_8.gated_control pin.t188 vss.t296 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X367 vdd.t307 PHI_1.t12 a_18728_1562# vdd.t306 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X368 vdd.t232 enable.t12 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t231 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X369 pin.t126 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 BUS[5].t13 vdd.t277 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X370 vdd.t7 a_3800_2002# a_3660_2122# vdd.t6 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X371 pin.t156 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 BUS[3].t9 vdd.t334 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X372 BUS[6].t3 swmatrix_Tgate_6.gated_control pin.t34 vss.t72 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X373 vss.t261 PHI_1.t13 a_6248_1562# vss.t260 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X374 pin.t3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[8].t0 vdd.t17 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X375 a_57004_1577# ShiftReg_row_10_2$1_0.Q[9] vss.t324 vss.t323 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X376 pin.t69 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[4].t6 vdd.t202 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X377 a_40896_2122# a_40380_1580# a_40748_1577# vss.t38 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X378 a_6716_1580# a_6248_1562# vdd.t41 vdd.t40 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X379 pin.t136 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 BUS[2].t3 vdd.t301 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X380 a_51256_2002# a_50912_2122# vss.t96 vss.t95 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X381 BUS[7].t10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t40 vdd.t73 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X382 a_7084_2122# ShiftReg_row_10_2$1_0.Q[1] vdd.t87 vdd.t86 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X383 vdd.t414 a_38776_2002# a_38636_2122# vdd.t413 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X384 pin.t108 swmatrix_Tgate_3.gated_control BUS[8].t5 vss.t209 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X385 pin.t33 swmatrix_Tgate_6.gated_control BUS[6].t2 vss.t71 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X386 a_47380_1577# a_46152_1562# a_47136_2122# vss.t55 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X387 a_16280_2002# a_15936_2122# vss.t339 vss.t338 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X388 BUS[6].t13 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t119 vdd.t252 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X389 a_476_1580# a_8_1562# vss.t61 vss.t60 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X390 BUS[4].t5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t178 vdd.t360 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X391 BUS[2].t9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t165 vdd.t347 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X392 BUS[1].t20 swmatrix_Tgate_9.gated_control pin.t96 vss.t199 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X393 vss.t267 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t266 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X394 swmatrix_Tgate_9.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t366 vss.t365 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X395 vdd.t526 PHI_2.t12 a_27432_1562# vdd.t525 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X396 BUS[10].t4 swmatrix_Tgate_2.gated_control pin.t15 vss.t25 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X397 vdd.t95 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] vdd.t94 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X398 a_53720_2002# a_53376_2122# vss.t368 vss.t367 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X399 vss.t403 PHI_2.t13 a_8712_1562# vss.t402 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X400 pin.t120 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[6].t12 vdd.t253 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X401 BUS[9].t11 swmatrix_Tgate_1.gated_control pin.t193 vss.t306 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X402 a_44524_2122# ShiftReg_row_10_2$1_0.Q[7] vdd.t451 vdd.t450 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X403 vss.t50 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss.t49 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X404 a_59616_2122# a_59100_1580# a_59468_1577# vss.t64 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X405 vdd.t234 enable.t13 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t233 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X406 vdd.t490 a_47480_2002# a_47340_2122# vdd.t489 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X407 pin.t223 swmatrix_Tgate_7.gated_control BUS[4].t19 vss.t385 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X408 a_51116_2122# a_50396_1580# a_50912_2122# vdd.t427 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X409 BUS[3].t8 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 pin.t170 vdd.t352 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X410 a_32044_1577# ShiftReg_row_10_2$1_0.Q[5] vss.t130 vss.t129 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X411 BUS[10].t13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t131 vdd.t296 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X412 pin.t55 swmatrix_Tgate_4.gated_control BUS[3].t20 vss.t101 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X413 vss.t121 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] vss.t120 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X414 a_36121_1539# ShiftReg_row_10_2$1_0.Q[6] vss.t174 vss.t173 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X415 BUS[7].t9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 pin.t39 vdd.t72 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X416 vdd.t182 a_20056_2002# a_19916_2122# vdd.t181 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X417 a_3456_2122# a_2940_1580# a_3308_1577# vss.t131 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X418 vdd.t59 a_13816_2002# a_13676_2122# vdd.t58 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X419 a_46988_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t27 vdd.t26 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X420 a_22420_1577# a_21192_1562# a_22176_2122# vss.t31 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X421 a_40896_2122# a_39912_1562# a_40748_2122# vdd.t367 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X422 pin.t161 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[10].t12 vdd.t343 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X423 pin.t179 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[4].t4 vdd.t361 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X424 vdd.t115 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t114 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X425 a_38432_2122# a_37916_1580# a_38284_1577# vss.t250 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X426 BUS[6].t11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t82 vdd.t215 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X427 BUS[2].t6 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 pin.t157 vdd.t337 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X428 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[9] vdd.t419 vdd.t418 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X429 BUS[4].t3 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 pin.t180 vdd.t362 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X430 vdd.t120 a_22520_2002# a_22380_2122# vdd.t119 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X431 vss.t263 PHI_1.t14 a_24968_1562# vss.t262 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X432 vss.t265 PHI_1.t15 a_18728_1562# vss.t264 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X433 a_59616_2122# a_58632_1562# a_59468_2122# vdd.t392 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X434 a_35000_2002# a_34656_2122# vdd.t144 vdd.t143 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X435 BUS[9].t10 swmatrix_Tgate_1.gated_control pin.t192 vss.t305 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X436 vss.t399 a_51256_2002# a_51156_1577# vss.t398 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X437 a_25436_1580# a_24968_1562# vdd.t515 vdd.t514 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X438 pin.t38 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 BUS[7].t8 vdd.t71 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X439 a_50396_1580# a_49928_1562# vss.t289 vss.t288 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X440 a_22028_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t170 vdd.t169 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X441 vss.t70 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t69 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X442 pin.t171 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 BUS[3].t7 vdd.t353 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X443 pin.t150 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 BUS[10].t11 vdd.t328 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X444 a_59468_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t303 vss.t302 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X445 a_32396_2122# a_31676_1580# a_32192_2122# vdd.t100 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X446 swmatrix_Tgate_7.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t40 vss.t39 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X447 swmatrix_Tgate_5.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t12 vdd.t11 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X448 BUS[9].t22 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t233 vdd.t529 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X449 a_3456_2122# a_2472_1562# a_3308_2122# vdd.t111 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X450 a_9548_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t150 vdd.t149 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X451 vss.t276 a_16280_2002# a_16180_1577# vss.t275 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X452 BUS[7].t7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t37 vdd.t70 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X453 pin.t54 swmatrix_Tgate_4.gated_control BUS[3].t19 vss.t100 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X454 swmatrix_Tgate_4.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t89 vss.t88 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X455 BUS[1].t7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 pin.t182 vdd.t389 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X456 a_15420_1580# a_14952_1562# vss.t229 vss.t228 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X457 vss.t328 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] vss.t327 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X458 BUS[5].t12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 pin.t237 vdd.t537 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X459 a_17401_1539# ShiftReg_row_10_2$1_0.Q[3] vss.t159 vss.t158 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X460 vss.t405 PHI_2.t14 a_27432_1562# vss.t404 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X461 a_844_1577# D_in.t1 vss.t246 vss.t245 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X462 a_3308_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t152 vss.t151 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X463 a_34140_1580# a_33672_1562# vdd.t323 vdd.t322 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X464 BUS[5].t1 swmatrix_Tgate_5.gated_control pin.t10 vss.t13 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X465 vss.t222 a_53720_2002# a_53620_1577# vss.t221 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X466 a_27900_1580# a_27432_1562# vdd.t482 vdd.t481 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X467 BUS[3].t18 swmatrix_Tgate_4.gated_control pin.t58 vss.t99 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X468 pin.t183 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 BUS[1].t6 vdd.t390 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X469 vdd.t241 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t240 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X470 pin.t238 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 BUS[5].t11 vdd.t538 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X471 a_52860_1580# a_52392_1562# vss.t189 vss.t188 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X472 a_38432_2122# a_37448_1562# a_38284_2122# vdd.t266 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X473 BUS[4].t18 swmatrix_Tgate_7.gated_control pin.t222 vss.t384 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X474 a_13816_2002# a_13472_2122# vdd.t410 vdd.t409 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X475 pin.t83 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[6].t10 vdd.t216 pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X476 a_50912_2122# a_50396_1580# a_50764_1577# vss.t331 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X477 a_34860_2122# a_34140_1580# a_34656_2122# vdd.t153 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X478 a_57396_1577# a_56168_1562# a_57152_2122# vss.t390 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X479 BUS[3].t6 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 pin.t129 vdd.t292 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X480 pin.t32 swmatrix_Tgate_6.gated_control BUS[6].t1 vss.t68 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X481 a_22176_2122# a_21660_1580# a_22028_1577# vss.t277 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X482 a_38284_1577# ShiftReg_row_10_2$1_0.Q[6] vss.t172 vss.t171 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X483 vss.t333 a_7576_2002# a_7476_1577# vss.t332 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X484 a_15936_2122# a_15420_1580# a_15788_1577# vss.t122 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X485 vdd.t273 PHI_1.t16 a_37448_1562# vdd.t272 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X486 BUS[8].t1 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t4 vdd.t18 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X487 a_51256_2002# a_50912_2122# vdd.t102 vdd.t101 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X488 vdd.t56 enable.t14 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t55 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X489 BUS[2].t7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 pin.t158 vdd.t338 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X490 vdd.t534 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t533 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X491 a_16280_2002# a_15936_2122# vdd.t435 vdd.t434 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X492 vdd.t497 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t496 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X493 pin.t184 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 BUS[1].t5 vdd.t391 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X494 pin.t239 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[5].t10 vdd.t539 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X495 pin.t172 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[2].t12 vdd.t354 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X496 pin.t95 swmatrix_Tgate_9.gated_control BUS[1].t19 vss.t198 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X497 vdd.t439 a_57496_2002# a_57356_2122# vdd.t438 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X498 a_59860_1577# a_58632_1562# a_59616_2122# vss.t291 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X499 a_35000_2002# a_34656_2122# vss.t141 vss.t140 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X500 BUS[1].t4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 pin.t229 vdd.t504 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X501 vss.t379 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] vss.t378 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X502 pin.t18 swmatrix_Tgate_2.gated_control BUS[10].t3 vss.t24 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X503 vss.t279 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t278 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X504 vdd.t528 PHI_2.t15 a_46152_1562# vdd.t527 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X505 a_32436_1577# a_31208_1562# a_32192_2122# vss.t137 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X506 BUS[6].t9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 pin.t84 vdd.t217 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X507 vdd.t364 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t363 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X508 BUS[10].t2 swmatrix_Tgate_2.gated_control pin.t17 vss.t23 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X509 a_3700_1577# a_2472_1562# a_3456_2122# vss.t109 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X510 a_13324_1577# ShiftReg_row_10_2$1_0.Q[2] vss.t349 vss.t348 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X511 pin.t137 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 BUS[3].t5 vdd.t302 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X512 a_57004_2122# ShiftReg_row_10_2$1_0.Q[9] vdd.t417 vdd.t416 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X513 a_50912_2122# a_49928_1562# a_50764_2122# vdd.t384 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X514 pin.t151 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[10].t10 vdd.t329 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X515 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t15 a_17401_1539# vss.t63 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X516 vdd.t1 enable.t16 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t0 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X517 pin.t210 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 BUS[8].t15 vdd.t467 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X518 pin.t74 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 BUS[6].t8 vdd.t207 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X519 vdd.t129 a_59960_2002# a_59820_2122# vdd.t128 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X520 a_28268_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t127 vdd.t126 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X521 a_22176_2122# a_21192_1562# a_22028_2122# vdd.t28 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X522 a_15936_2122# a_14952_1562# a_15788_2122# vdd.t269 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X523 a_50764_1577# ShiftReg_row_10_2$1_0.Q[8] vss.t166 vss.t165 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X524 pin.t190 swmatrix_Tgate_8.gated_control BUS[2].t17 vss.t295 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X525 BUS[10].t9 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 pin.t148 vdd.t326 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X526 BUS[1].t3 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 pin.t230 vdd.t505 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X527 BUS[8].t16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 pin.t211 vdd.t468 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X528 vdd.t176 a_32536_2002# a_32396_2122# vdd.t175 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X529 BUS[4].t2 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t72 vdd.t205 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X530 a_13816_2002# a_13472_2122# vss.t319 vss.t318 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X531 a_41140_1577# a_39912_1562# a_40896_2122# vss.t270 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X532 a_15788_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t274 vss.t273 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X533 a_10040_2002# a_9696_2122# vss.t85 vss.t84 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X534 BUS[9].t23 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 pin.t234 vdd.t530 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X535 BUS[7].t6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 pin.t36 vdd.t69 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X536 vdd.t122 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] vdd.t121 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X537 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[6] vdd.t178 vdd.t177 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X538 pin.t231 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 BUS[1].t2 vdd.t506 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X539 vdd.t520 PHI_2.t16 a_21192_1562# vdd.t519 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X540 pin.t173 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 BUS[2].t13 vdd.t355 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X541 vss.t178 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] vss.t177 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X542 pin.t128 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 BUS[9].t1 vdd.t291 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X543 a_57152_2122# a_56636_1580# a_57004_1577# vss.t322 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X544 vss.t372 a_26296_2002# a_26196_1577# vss.t371 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X545 BUS[2].t1 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t134 vdd.t299 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X546 pin.t191 swmatrix_Tgate_1.gated_control BUS[9].t9 vss.t304 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X547 vdd.t158 a_41240_2002# a_41100_2122# vdd.t157 pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X548 a_25436_1580# a_24968_1562# vss.t396 vss.t395 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X549 BUS[8].t17 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t212 vdd.t477 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X550 vss.t232 PHI_1.t17 a_37448_1562# vss.t231 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X551 a_13716_1577# a_12488_1562# a_13472_2122# vss.t75 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X552 BUS[3].t4 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 pin.t138 vdd.t303 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X553 a_44156_1580# a_43688_1562# vdd.t193 vdd.t192 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X554 a_37916_1580# a_37448_1562# vdd.t265 vdd.t264 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X555 pin.t149 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 BUS[10].t8 vdd.t327 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X556 BUS[1].t18 swmatrix_Tgate_9.gated_control pin.t94 vss.t197 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X557 pin.t213 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[8].t18 vdd.t478 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X558 a_40748_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t110 vdd.t109 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X559 pin.t91 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 BUS[5].t9 vdd.t226 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X560 pin.t35 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[7].t13 vdd.t68 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X561 a_44876_2122# a_44156_1580# a_44672_2122# vdd.t44 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X562 vss.t351 a_35000_2002# a_34900_1577# vss.t350 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X563 vss.t91 a_28760_2002# a_28660_1577# vss.t90 nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X564 swmatrix_Tgate_6.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t59 vss.t58 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X565 swmatrix_Tgate_0.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t268 vdd.t267 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X566 vss.t208 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t207 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X567 a_34140_1580# a_33672_1562# vss.t256 vss.t255 nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X568 BUS[4].t1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 pin.t73 vdd.t206 pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X569 a_29881_1539# ShiftReg_row_10_2$1_0.Q[5] vss.t128 vss.t127 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X570 vss.t401 PHI_2.t17 a_46152_1562# vss.t400 nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X571 a_992_2122# a_476_1580# a_844_1577# vss.t20 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X572 BUS[9].t2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t141 vdd.t310 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X573 a_46620_1580# a_46152_1562# vdd.t48 vdd.t47 pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X574 a_7576_2002# a_7232_2122# vss.t343 vss.t342 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X575 a_16140_2122# a_15420_1580# a_15936_2122# vdd.t125 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X576 vdd.t426 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] vdd.t425 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X577 pin.t139 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[2].t4 vdd.t308 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X578 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN ShiftReg_row_10_2$1_0.Q[3] vdd.t165 vdd.t164 pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X579 vss.t317 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t316 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X580 vdd.t25 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t24 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X581 BUS[7].t1 swmatrix_Tgate_0.gated_control pin.t21 vss.t48 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X582 a_57152_2122# a_56168_1562# a_57004_2122# vdd.t499 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X583 BUS[5].t0 swmatrix_Tgate_5.gated_control pin.t9 vss.t12 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X584 a_26296_2002# a_25952_2122# vdd.t456 vdd.t455 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X585 pin.t142 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[9].t3 vdd.t311 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X586 a_53580_2122# a_52860_1580# a_53376_2122# vdd.t315 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X587 pin.t103 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 BUS[3].t3 vdd.t238 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X588 pin.t147 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[10].t7 vdd.t325 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X589 vss.t383 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss.t382 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X590 vss.t94 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t93 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X591 a_34656_2122# a_34140_1580# a_34508_1577# vss.t150 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X592 pin.t20 swmatrix_Tgate_0.gated_control BUS[7].t0 vss.t47 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X593 vdd.t275 PHI_1.t18 a_56168_1562# vdd.t274 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X594 a_53228_1577# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss.t98 vss.t97 nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X595 BUS[5].t8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t92 vdd.t227 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X596 BUS[3].t2 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 pin.t104 vdd.t239 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X597 a_3308_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t156 vdd.t155 pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X598 BUS[10].t6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 pin.t146 vdd.t324 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X599 swmatrix_Tgate_8.gated_control ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss.t216 vss.t215 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X600 vss.t362 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] vss.t361 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X601 a_28760_2002# a_28416_2122# vdd.t424 vdd.t423 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X602 a_7436_2122# a_6716_1580# a_7232_2122# vdd.t454 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X603 a_11161_1539# ShiftReg_row_10_2$1_0.Q[2] vss.t347 vss.t346 nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
X604 vss.t337 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] vss.t336 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X605 BUS[2].t5 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 pin.t140 vdd.t309 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X606 vdd.t396 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t395 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X607 vdd.t230 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t229 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X608 pin.t70 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[1].t1 vdd.t203 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X609 BUS[10].t1 swmatrix_Tgate_2.gated_control pin.t14 vss.t22 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X610 pin.t93 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[5].t7 vdd.t228 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X611 pin.t201 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[9].t15 vdd.t420 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X612 pin.t75 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 BUS[6].t7 vdd.t208 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X613 pin.t117 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[4].t0 vdd.t250 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X614 vss.t133 a_59616_2122# d_out.t0 vss.t132 nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X615 a_47480_2002# a_47136_2122# vss.t119 vss.t118 nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X616 a_992_2122# a_8_1562# a_844_2122# vdd.t52 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X617 pin.t13 swmatrix_Tgate_2.gated_control BUS[10].t0 vss.t21 nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X618 vdd.t522 PHI_2.t18 a_58632_1562# vdd.t521 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X619 a_51156_1577# a_49928_1562# a_50912_2122# vss.t287 nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X620 vdd.t493 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] vdd.t492 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X621 a_13472_2122# a_12956_1580# a_13324_1577# vss.t183 nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X622 BUS[6].t6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 pin.t181 vdd.t388 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X623 BUS[3].t1 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 pin.t76 vdd.t209 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X624 vdd.t376 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd.t375 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X625 vdd.t336 PHI_1.t19 a_31208_1562# vdd.t335 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X626 a_9900_2122# a_9180_1580# a_9696_2122# vdd.t148 pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
X627 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t17 a_36121_1539# vss.t0 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X628 vdd.t3 enable.t18 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd.t2 pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X629 BUS[2].t16 swmatrix_Tgate_8.gated_control pin.t189 vss.t294 nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X630 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable.t19 a_29881_1539# vss.t1 nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X631 pin.t71 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[1].t0 vdd.t204 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X632 vdd.t524 PHI_2.t19 a_2472_1562# vdd.t523 pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X633 pin.t216 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[8].t19 vdd.t484 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X634 pin.t90 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[5].t6 vdd.t225 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X635 vdd.t400 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vdd.t399 pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X636 pin.t232 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 BUS[3].t0 vdd.t507 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X637 a_10040_2002# a_9696_2122# vdd.t93 vdd.t92 pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X638 a_34656_2122# a_33672_1562# a_34508_2122# vdd.t321 pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X639 BUS[6].t0 swmatrix_Tgate_6.gated_control pin.t31 vss.t67 nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
R0 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.7994
R1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R3 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R4 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R8 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R13 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R17 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R18 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R19 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 4.63372
R20 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 3.85252
R21 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R22 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R23 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R24 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R25 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R26 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R27 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R28 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R29 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R30 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R31 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R32 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R33 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R34 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R35 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R36 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R37 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R38 BUS[7].n2 BUS[7].n0 15.3751
R39 BUS[7].n9 BUS[7].n7 15.2168
R40 BUS[7].n2 BUS[7].n1 15.0151
R41 BUS[7].n4 BUS[7].n3 15.0151
R42 BUS[7].n21 BUS[7].n20 14.8568
R43 BUS[7].n19 BUS[7].n18 14.8568
R44 BUS[7].n17 BUS[7].n16 14.8568
R45 BUS[7].n15 BUS[7].n14 14.8568
R46 BUS[7].n13 BUS[7].n12 14.8568
R47 BUS[7].n11 BUS[7].n10 14.8568
R48 BUS[7].n9 BUS[7].n8 14.8568
R49 BUS[7].n6 BUS[7].n5 14.8568
R50 BUS[7].n22 BUS[7] 0.921051
R51 BUS[7].n6 BUS[7].n4 0.8825
R52 BUS[7].n20 BUS[7].t22 0.4555
R53 BUS[7].n20 BUS[7].t10 0.4555
R54 BUS[7].n18 BUS[7].t8 0.4555
R55 BUS[7].n18 BUS[7].t11 0.4555
R56 BUS[7].n16 BUS[7].t20 0.4555
R57 BUS[7].n16 BUS[7].t21 0.4555
R58 BUS[7].n14 BUS[7].t13 0.4555
R59 BUS[7].n14 BUS[7].t7 0.4555
R60 BUS[7].n12 BUS[7].t17 0.4555
R61 BUS[7].n12 BUS[7].t14 0.4555
R62 BUS[7].n10 BUS[7].t23 0.4555
R63 BUS[7].n10 BUS[7].t9 0.4555
R64 BUS[7].n8 BUS[7].t19 0.4555
R65 BUS[7].n8 BUS[7].t12 0.4555
R66 BUS[7].n7 BUS[7].t16 0.4555
R67 BUS[7].n7 BUS[7].t6 0.4555
R68 BUS[7].n5 BUS[7].t18 0.4555
R69 BUS[7].n5 BUS[7].t15 0.4555
R70 BUS[7].n0 BUS[7].t3 0.41
R71 BUS[7].n0 BUS[7].t1 0.41
R72 BUS[7].n1 BUS[7].t0 0.41
R73 BUS[7].n1 BUS[7].t2 0.41
R74 BUS[7].n3 BUS[7].t4 0.41
R75 BUS[7].n3 BUS[7].t5 0.41
R76 BUS[7].n4 BUS[7].n2 0.3605
R77 BUS[7].n11 BUS[7].n9 0.3605
R78 BUS[7].n13 BUS[7].n11 0.3605
R79 BUS[7].n15 BUS[7].n13 0.3605
R80 BUS[7].n17 BUS[7].n15 0.3605
R81 BUS[7].n19 BUS[7].n17 0.3605
R82 BUS[7].n21 BUS[7].n19 0.3605
R83 BUS[7].n22 BUS[7].n6 0.203
R84 BUS[7] BUS[7].n22 0.0430197
R85 BUS[7].n22 BUS[7].n21 0.015125
R86 pin.n100 pin.t150 11.5218
R87 pin.n109 pin.t13 11.3429
R88 pin.n112 pin.t15 11.3429
R89 pin.n123 pin.t195 11.3429
R90 pin.n126 pin.t192 11.3429
R91 pin.n137 pin.t109 11.3429
R92 pin.n140 pin.t106 11.3429
R93 pin.n151 pin.t24 11.3429
R94 pin.n154 pin.t21 11.3429
R95 pin.n165 pin.t33 11.3429
R96 pin.n168 pin.t31 11.3429
R97 pin.n179 pin.t7 11.3429
R98 pin.n182 pin.t10 11.3429
R99 pin.n193 pin.t227 11.3429
R100 pin.n196 pin.t226 11.3429
R101 pin.n207 pin.t55 11.3429
R102 pin.n210 pin.t57 11.3429
R103 pin.n221 pin.t187 11.3429
R104 pin.n224 pin.t186 11.3429
R105 pin.n235 pin.t98 11.3429
R106 pin.n238 pin.t96 11.3429
R107 pin.n108 pin.t200 11.2918
R108 pin.n113 pin.t204 11.2918
R109 pin.n122 pin.t168 11.2918
R110 pin.n127 pin.t217 11.2918
R111 pin.n136 pin.t209 11.2918
R112 pin.n141 pin.t52 11.2918
R113 pin.n150 pin.t51 11.2918
R114 pin.n155 pin.t83 11.2918
R115 pin.n164 pin.t122 11.2918
R116 pin.n169 pin.t238 11.2918
R117 pin.n178 pin.t125 11.2918
R118 pin.n183 pin.t68 11.2918
R119 pin.n192 pin.t73 11.2918
R120 pin.n197 pin.t64 11.2918
R121 pin.n206 pin.t170 11.2918
R122 pin.n211 pin.t219 11.2918
R123 pin.n220 pin.t167 11.2918
R124 pin.n225 pin.t183 11.2918
R125 pin.n234 pin.t230 11.2918
R126 pin.n110 pin.n91 10.7129
R127 pin.n111 pin.n90 10.7129
R128 pin.n124 pin.n81 10.7129
R129 pin.n125 pin.n80 10.7129
R130 pin.n138 pin.n71 10.7129
R131 pin.n139 pin.n70 10.7129
R132 pin.n152 pin.n61 10.7129
R133 pin.n153 pin.n60 10.7129
R134 pin.n166 pin.n51 10.7129
R135 pin.n167 pin.n50 10.7129
R136 pin.n180 pin.n41 10.7129
R137 pin.n181 pin.n40 10.7129
R138 pin.n194 pin.n31 10.7129
R139 pin.n195 pin.n30 10.7129
R140 pin.n208 pin.n21 10.7129
R141 pin.n209 pin.n20 10.7129
R142 pin.n222 pin.n11 10.7129
R143 pin.n223 pin.n10 10.7129
R144 pin.n236 pin.n1 10.7129
R145 pin.n237 pin.n0 10.7129
R146 pin.n100 pin.n99 10.5568
R147 pin.n101 pin.n98 10.5568
R148 pin.n102 pin.n97 10.5568
R149 pin.n103 pin.n96 10.5568
R150 pin.n104 pin.n95 10.5568
R151 pin.n105 pin.n94 10.5568
R152 pin.n106 pin.n93 10.5568
R153 pin.n107 pin.n92 10.5568
R154 pin.n114 pin.n89 10.5568
R155 pin.n115 pin.n88 10.5568
R156 pin.n116 pin.n87 10.5568
R157 pin.n117 pin.n86 10.5568
R158 pin.n118 pin.n85 10.5568
R159 pin.n119 pin.n84 10.5568
R160 pin.n120 pin.n83 10.5568
R161 pin.n121 pin.n82 10.5568
R162 pin.n128 pin.n79 10.5568
R163 pin.n129 pin.n78 10.5568
R164 pin.n130 pin.n77 10.5568
R165 pin.n131 pin.n76 10.5568
R166 pin.n132 pin.n75 10.5568
R167 pin.n133 pin.n74 10.5568
R168 pin.n134 pin.n73 10.5568
R169 pin.n135 pin.n72 10.5568
R170 pin.n142 pin.n69 10.5568
R171 pin.n143 pin.n68 10.5568
R172 pin.n144 pin.n67 10.5568
R173 pin.n145 pin.n66 10.5568
R174 pin.n146 pin.n65 10.5568
R175 pin.n147 pin.n64 10.5568
R176 pin.n148 pin.n63 10.5568
R177 pin.n149 pin.n62 10.5568
R178 pin.n156 pin.n59 10.5568
R179 pin.n157 pin.n58 10.5568
R180 pin.n158 pin.n57 10.5568
R181 pin.n159 pin.n56 10.5568
R182 pin.n160 pin.n55 10.5568
R183 pin.n161 pin.n54 10.5568
R184 pin.n162 pin.n53 10.5568
R185 pin.n163 pin.n52 10.5568
R186 pin.n170 pin.n49 10.5568
R187 pin.n171 pin.n48 10.5568
R188 pin.n172 pin.n47 10.5568
R189 pin.n173 pin.n46 10.5568
R190 pin.n174 pin.n45 10.5568
R191 pin.n175 pin.n44 10.5568
R192 pin.n176 pin.n43 10.5568
R193 pin.n177 pin.n42 10.5568
R194 pin.n184 pin.n39 10.5568
R195 pin.n185 pin.n38 10.5568
R196 pin.n186 pin.n37 10.5568
R197 pin.n187 pin.n36 10.5568
R198 pin.n188 pin.n35 10.5568
R199 pin.n189 pin.n34 10.5568
R200 pin.n190 pin.n33 10.5568
R201 pin.n191 pin.n32 10.5568
R202 pin.n198 pin.n29 10.5568
R203 pin.n199 pin.n28 10.5568
R204 pin.n200 pin.n27 10.5568
R205 pin.n201 pin.n26 10.5568
R206 pin.n202 pin.n25 10.5568
R207 pin.n203 pin.n24 10.5568
R208 pin.n204 pin.n23 10.5568
R209 pin.n205 pin.n22 10.5568
R210 pin.n212 pin.n19 10.5568
R211 pin.n213 pin.n18 10.5568
R212 pin.n214 pin.n17 10.5568
R213 pin.n215 pin.n16 10.5568
R214 pin.n216 pin.n15 10.5568
R215 pin.n217 pin.n14 10.5568
R216 pin.n218 pin.n13 10.5568
R217 pin.n219 pin.n12 10.5568
R218 pin.n226 pin.n9 10.5568
R219 pin.n227 pin.n8 10.5568
R220 pin.n228 pin.n7 10.5568
R221 pin.n229 pin.n6 10.5568
R222 pin.n230 pin.n5 10.5568
R223 pin.n231 pin.n4 10.5568
R224 pin.n232 pin.n3 10.5568
R225 pin.n233 pin.n2 10.5568
R226 pin.n225 pin 0.99904
R227 pin.n113 pin 0.67123
R228 pin.n127 pin 0.67123
R229 pin.n141 pin 0.67123
R230 pin.n155 pin 0.67123
R231 pin.n169 pin 0.67123
R232 pin.n183 pin 0.67123
R233 pin.n197 pin 0.67123
R234 pin.n211 pin 0.67123
R235 pin pin.n112 0.564807
R236 pin pin.n126 0.564807
R237 pin pin.n140 0.564807
R238 pin pin.n154 0.564807
R239 pin pin.n168 0.564807
R240 pin pin.n182 0.564807
R241 pin pin.n196 0.564807
R242 pin pin.n210 0.564807
R243 pin pin.n224 0.564807
R244 pin pin.n238 0.564807
R245 pin.n99 pin.t130 0.4555
R246 pin.n99 pin.t228 0.4555
R247 pin.n98 pin.t146 0.4555
R248 pin.n98 pin.t163 0.4555
R249 pin.n97 pin.t77 0.4555
R250 pin.n97 pin.t147 0.4555
R251 pin.n96 pin.t78 0.4555
R252 pin.n96 pin.t132 0.4555
R253 pin.n95 pin.t148 0.4555
R254 pin.n95 pin.t161 0.4555
R255 pin.n94 pin.t164 0.4555
R256 pin.n94 pin.t151 0.4555
R257 pin.n93 pin.t131 0.4555
R258 pin.n93 pin.t162 0.4555
R259 pin.n92 pin.t133 0.4555
R260 pin.n92 pin.t149 0.4555
R261 pin.n89 pin.t59 0.4555
R262 pin.n89 pin.t128 0.4555
R263 pin.n88 pin.t215 0.4555
R264 pin.n88 pin.t177 0.4555
R265 pin.n87 pin.t234 0.4555
R266 pin.n87 pin.t142 0.4555
R267 pin.n86 pin.t160 0.4555
R268 pin.n86 pin.t202 0.4555
R269 pin.n85 pin.t141 0.4555
R270 pin.n85 pin.t205 0.4555
R271 pin.n84 pin.t214 0.4555
R272 pin.n84 pin.t176 0.4555
R273 pin.n83 pin.t233 0.4555
R274 pin.n83 pin.t169 0.4555
R275 pin.n82 pin.t203 0.4555
R276 pin.n82 pin.t201 0.4555
R277 pin.n79 pin.t4 0.4555
R278 pin.n79 pin.t3 0.4555
R279 pin.n78 pin.t236 0.4555
R280 pin.n78 pin.t216 0.4555
R281 pin.n77 pin.t211 0.4555
R282 pin.n77 pin.t206 0.4555
R283 pin.n76 pin.t5 0.4555
R284 pin.n76 pin.t210 0.4555
R285 pin.n75 pin.t6 0.4555
R286 pin.n75 pin.t218 0.4555
R287 pin.n74 pin.t235 0.4555
R288 pin.n74 pin.t213 0.4555
R289 pin.n73 pin.t208 0.4555
R290 pin.n73 pin.t19 0.4555
R291 pin.n72 pin.t212 0.4555
R292 pin.n72 pin.t207 0.4555
R293 pin.n69 pin.t36 0.4555
R294 pin.n69 pin.t45 0.4555
R295 pin.n68 pin.t42 0.4555
R296 pin.n68 pin.t49 0.4555
R297 pin.n67 pin.t39 0.4555
R298 pin.n67 pin.t43 0.4555
R299 pin.n66 pin.t50 0.4555
R300 pin.n66 pin.t35 0.4555
R301 pin.n65 pin.t37 0.4555
R302 pin.n65 pin.t46 0.4555
R303 pin.n64 pin.t47 0.4555
R304 pin.n64 pin.t38 0.4555
R305 pin.n63 pin.t41 0.4555
R306 pin.n63 pin.t48 0.4555
R307 pin.n62 pin.t40 0.4555
R308 pin.n62 pin.t44 0.4555
R309 pin.n59 pin.t118 0.4555
R310 pin.n59 pin.t87 0.4555
R311 pin.n58 pin.t181 0.4555
R312 pin.n58 pin.t74 0.4555
R313 pin.n57 pin.t86 0.4555
R314 pin.n57 pin.t75 0.4555
R315 pin.n56 pin.t84 0.4555
R316 pin.n56 pin.t120 0.4555
R317 pin.n55 pin.t89 0.4555
R318 pin.n55 pin.t121 0.4555
R319 pin.n54 pin.t119 0.4555
R320 pin.n54 pin.t88 0.4555
R321 pin.n53 pin.t102 0.4555
R322 pin.n53 pin.t123 0.4555
R323 pin.n52 pin.t82 0.4555
R324 pin.n52 pin.t85 0.4555
R325 pin.n49 pin.t1 0.4555
R326 pin.n49 pin.t91 0.4555
R327 pin.n48 pin.t237 0.4555
R328 pin.n48 pin.t0 0.4555
R329 pin.n47 pin.t100 0.4555
R330 pin.n47 pin.t93 0.4555
R331 pin.n46 pin.t28 0.4555
R332 pin.n46 pin.t26 0.4555
R333 pin.n45 pin.t92 0.4555
R334 pin.n45 pin.t239 0.4555
R335 pin.n44 pin.t2 0.4555
R336 pin.n44 pin.t101 0.4555
R337 pin.n43 pin.t154 0.4555
R338 pin.n43 pin.t126 0.4555
R339 pin.n42 pin.t27 0.4555
R340 pin.n42 pin.t90 0.4555
R341 pin.n39 pin.t66 0.4555
R342 pin.n39 pin.t117 0.4555
R343 pin.n38 pin.t67 0.4555
R344 pin.n38 pin.t65 0.4555
R345 pin.n37 pin.t114 0.4555
R346 pin.n37 pin.t79 0.4555
R347 pin.n36 pin.t178 0.4555
R348 pin.n36 pin.t81 0.4555
R349 pin.n35 pin.t60 0.4555
R350 pin.n35 pin.t69 0.4555
R351 pin.n34 pin.t180 0.4555
R352 pin.n34 pin.t116 0.4555
R353 pin.n33 pin.t72 0.4555
R354 pin.n33 pin.t179 0.4555
R355 pin.n32 pin.t115 0.4555
R356 pin.n32 pin.t80 0.4555
R357 pin.n29 pin.t138 0.4555
R358 pin.n29 pin.t171 0.4555
R359 pin.n28 pin.t199 0.4555
R360 pin.n28 pin.t127 0.4555
R361 pin.n27 pin.t104 0.4555
R362 pin.n27 pin.t62 0.4555
R363 pin.n26 pin.t61 0.4555
R364 pin.n26 pin.t103 0.4555
R365 pin.n25 pin.t129 0.4555
R366 pin.n25 pin.t156 0.4555
R367 pin.n24 pin.t63 0.4555
R368 pin.n24 pin.t232 0.4555
R369 pin.n23 pin.t155 0.4555
R370 pin.n23 pin.t221 0.4555
R371 pin.n22 pin.t76 0.4555
R372 pin.n22 pin.t137 0.4555
R373 pin.n19 pin.t140 0.4555
R374 pin.n19 pin.t172 0.4555
R375 pin.n18 pin.t165 0.4555
R376 pin.n18 pin.t174 0.4555
R377 pin.n17 pin.t158 0.4555
R378 pin.n17 pin.t136 0.4555
R379 pin.n16 pin.t220 0.4555
R380 pin.n16 pin.t124 0.4555
R381 pin.n15 pin.t134 0.4555
R382 pin.n15 pin.t166 0.4555
R383 pin.n14 pin.t175 0.4555
R384 pin.n14 pin.t173 0.4555
R385 pin.n13 pin.t157 0.4555
R386 pin.n13 pin.t135 0.4555
R387 pin.n12 pin.t159 0.4555
R388 pin.n12 pin.t139 0.4555
R389 pin.n9 pin.t113 0.4555
R390 pin.n9 pin.t111 0.4555
R391 pin.n8 pin.t182 0.4555
R392 pin.n8 pin.t153 0.4555
R393 pin.n7 pin.t198 0.4555
R394 pin.n7 pin.t70 0.4555
R395 pin.n6 pin.t229 0.4555
R396 pin.n6 pin.t144 0.4555
R397 pin.n5 pin.t112 0.4555
R398 pin.n5 pin.t184 0.4555
R399 pin.n4 pin.t143 0.4555
R400 pin.n4 pin.t152 0.4555
R401 pin.n3 pin.t197 0.4555
R402 pin.n3 pin.t231 0.4555
R403 pin.n2 pin.t145 0.4555
R404 pin.n2 pin.t71 0.4555
R405 pin.n91 pin.t17 0.41
R406 pin.n91 pin.t16 0.41
R407 pin.n90 pin.t14 0.41
R408 pin.n90 pin.t18 0.41
R409 pin.n81 pin.t193 0.41
R410 pin.n81 pin.t194 0.41
R411 pin.n80 pin.t196 0.41
R412 pin.n80 pin.t191 0.41
R413 pin.n71 pin.t110 0.41
R414 pin.n71 pin.t105 0.41
R415 pin.n70 pin.t107 0.41
R416 pin.n70 pin.t108 0.41
R417 pin.n61 pin.t25 0.41
R418 pin.n61 pin.t20 0.41
R419 pin.n60 pin.t22 0.41
R420 pin.n60 pin.t23 0.41
R421 pin.n51 pin.t29 0.41
R422 pin.n51 pin.t32 0.41
R423 pin.n50 pin.t34 0.41
R424 pin.n50 pin.t30 0.41
R425 pin.n41 pin.t9 0.41
R426 pin.n41 pin.t11 0.41
R427 pin.n40 pin.t8 0.41
R428 pin.n40 pin.t12 0.41
R429 pin.n31 pin.t222 0.41
R430 pin.n31 pin.t225 0.41
R431 pin.n30 pin.t224 0.41
R432 pin.n30 pin.t223 0.41
R433 pin.n21 pin.t58 0.41
R434 pin.n21 pin.t56 0.41
R435 pin.n20 pin.t53 0.41
R436 pin.n20 pin.t54 0.41
R437 pin.n11 pin.t188 0.41
R438 pin.n11 pin.t185 0.41
R439 pin.n10 pin.t189 0.41
R440 pin.n10 pin.t190 0.41
R441 pin.n1 pin.t94 0.41
R442 pin.n1 pin.t97 0.41
R443 pin.n0 pin.t99 0.41
R444 pin.n0 pin.t95 0.41
R445 pin.n109 pin.n108 0.266558
R446 pin.n123 pin.n122 0.266558
R447 pin.n137 pin.n136 0.266558
R448 pin.n151 pin.n150 0.266558
R449 pin.n165 pin.n164 0.266558
R450 pin.n179 pin.n178 0.266558
R451 pin.n193 pin.n192 0.266558
R452 pin.n207 pin.n206 0.266558
R453 pin.n221 pin.n220 0.266558
R454 pin.n235 pin.n234 0.266558
R455 pin.n108 pin.n107 0.230427
R456 pin.n114 pin.n113 0.230427
R457 pin.n122 pin.n121 0.230427
R458 pin.n128 pin.n127 0.230427
R459 pin.n136 pin.n135 0.230427
R460 pin.n142 pin.n141 0.230427
R461 pin.n150 pin.n149 0.230427
R462 pin.n156 pin.n155 0.230427
R463 pin.n164 pin.n163 0.230427
R464 pin.n170 pin.n169 0.230427
R465 pin.n178 pin.n177 0.230427
R466 pin.n184 pin.n183 0.230427
R467 pin.n192 pin.n191 0.230427
R468 pin.n198 pin.n197 0.230427
R469 pin.n206 pin.n205 0.230427
R470 pin.n212 pin.n211 0.230427
R471 pin.n220 pin.n219 0.230427
R472 pin.n226 pin.n225 0.230427
R473 pin.n234 pin.n233 0.230427
R474 pin.n110 pin.n109 0.22977
R475 pin.n124 pin.n123 0.22977
R476 pin.n138 pin.n137 0.22977
R477 pin.n152 pin.n151 0.22977
R478 pin.n166 pin.n165 0.22977
R479 pin.n180 pin.n179 0.22977
R480 pin.n194 pin.n193 0.22977
R481 pin.n208 pin.n207 0.22977
R482 pin.n222 pin.n221 0.22977
R483 pin.n236 pin.n235 0.22977
R484 pin.n112 pin.n111 0.227799
R485 pin.n126 pin.n125 0.227799
R486 pin.n140 pin.n139 0.227799
R487 pin.n154 pin.n153 0.227799
R488 pin.n168 pin.n167 0.227799
R489 pin.n182 pin.n181 0.227799
R490 pin.n196 pin.n195 0.227799
R491 pin.n210 pin.n209 0.227799
R492 pin.n224 pin.n223 0.227799
R493 pin.n238 pin.n237 0.227799
R494 pin.n101 pin.n100 0.210719
R495 pin.n102 pin.n101 0.210719
R496 pin.n103 pin.n102 0.210719
R497 pin.n104 pin.n103 0.210719
R498 pin.n105 pin.n104 0.210719
R499 pin.n106 pin.n105 0.210719
R500 pin.n107 pin.n106 0.210719
R501 pin.n111 pin.n110 0.210719
R502 pin.n115 pin.n114 0.210719
R503 pin.n116 pin.n115 0.210719
R504 pin.n117 pin.n116 0.210719
R505 pin.n118 pin.n117 0.210719
R506 pin.n119 pin.n118 0.210719
R507 pin.n120 pin.n119 0.210719
R508 pin.n121 pin.n120 0.210719
R509 pin.n125 pin.n124 0.210719
R510 pin.n129 pin.n128 0.210719
R511 pin.n130 pin.n129 0.210719
R512 pin.n131 pin.n130 0.210719
R513 pin.n132 pin.n131 0.210719
R514 pin.n133 pin.n132 0.210719
R515 pin.n134 pin.n133 0.210719
R516 pin.n135 pin.n134 0.210719
R517 pin.n139 pin.n138 0.210719
R518 pin.n143 pin.n142 0.210719
R519 pin.n144 pin.n143 0.210719
R520 pin.n145 pin.n144 0.210719
R521 pin.n146 pin.n145 0.210719
R522 pin.n147 pin.n146 0.210719
R523 pin.n148 pin.n147 0.210719
R524 pin.n149 pin.n148 0.210719
R525 pin.n153 pin.n152 0.210719
R526 pin.n157 pin.n156 0.210719
R527 pin.n158 pin.n157 0.210719
R528 pin.n159 pin.n158 0.210719
R529 pin.n160 pin.n159 0.210719
R530 pin.n161 pin.n160 0.210719
R531 pin.n162 pin.n161 0.210719
R532 pin.n163 pin.n162 0.210719
R533 pin.n167 pin.n166 0.210719
R534 pin.n171 pin.n170 0.210719
R535 pin.n172 pin.n171 0.210719
R536 pin.n173 pin.n172 0.210719
R537 pin.n174 pin.n173 0.210719
R538 pin.n175 pin.n174 0.210719
R539 pin.n176 pin.n175 0.210719
R540 pin.n177 pin.n176 0.210719
R541 pin.n181 pin.n180 0.210719
R542 pin.n185 pin.n184 0.210719
R543 pin.n186 pin.n185 0.210719
R544 pin.n187 pin.n186 0.210719
R545 pin.n188 pin.n187 0.210719
R546 pin.n189 pin.n188 0.210719
R547 pin.n190 pin.n189 0.210719
R548 pin.n191 pin.n190 0.210719
R549 pin.n195 pin.n194 0.210719
R550 pin.n199 pin.n198 0.210719
R551 pin.n200 pin.n199 0.210719
R552 pin.n201 pin.n200 0.210719
R553 pin.n202 pin.n201 0.210719
R554 pin.n203 pin.n202 0.210719
R555 pin.n204 pin.n203 0.210719
R556 pin.n205 pin.n204 0.210719
R557 pin.n209 pin.n208 0.210719
R558 pin.n213 pin.n212 0.210719
R559 pin.n214 pin.n213 0.210719
R560 pin.n215 pin.n214 0.210719
R561 pin.n216 pin.n215 0.210719
R562 pin.n217 pin.n216 0.210719
R563 pin.n218 pin.n217 0.210719
R564 pin.n219 pin.n218 0.210719
R565 pin.n223 pin.n222 0.210719
R566 pin.n227 pin.n226 0.210719
R567 pin.n228 pin.n227 0.210719
R568 pin.n229 pin.n228 0.210719
R569 pin.n230 pin.n229 0.210719
R570 pin.n231 pin.n230 0.210719
R571 pin.n232 pin.n231 0.210719
R572 pin.n233 pin.n232 0.210719
R573 pin.n237 pin.n236 0.210719
R574 vdd.t137 vdd.t135 667.707
R575 vdd.t375 vdd.t377 667.707
R576 vdd.t473 vdd.t471 667.707
R577 vdd.t103 vdd.t101 667.707
R578 vdd.t121 vdd.t123 667.707
R579 vdd.t13 vdd.t15 667.707
R580 vdd.t492 vdd.t494 667.707
R581 vdd.t363 vdd.t365 667.707
R582 vdd.t145 vdd.t143 667.707
R583 vdd.t319 vdd.t317 667.707
R584 vdd.t425 vdd.t423 667.707
R585 vdd.t457 vdd.t455 667.707
R586 vdd.t461 vdd.t459 667.707
R587 vdd.t533 vdd.t535 667.707
R588 vdd.t436 vdd.t434 667.707
R589 vdd.t411 vdd.t409 667.707
R590 vdd.t94 vdd.t92 667.707
R591 vdd.t440 vdd.t442 667.707
R592 vdd.t185 vdd.t183 667.707
R593 vdd.t114 vdd.t116 667.707
R594 vdd.n68 vdd.t229 652.42
R595 vdd.n71 vdd.t395 652.42
R596 vdd.n74 vdd.t107 652.42
R597 vdd.n77 vdd.t496 652.42
R598 vdd.n80 vdd.t21 652.42
R599 vdd.n83 vdd.t63 652.42
R600 vdd.n86 vdd.t45 652.42
R601 vdd.n89 vdd.t240 652.42
R602 vdd.n92 vdd.t399 652.42
R603 vdd.n95 vdd.t24 652.42
R604 vdd.t397 vdd.t393 574.104
R605 vdd.t416 vdd.t500 574.104
R606 vdd.t105 vdd.t195 574.104
R607 vdd.t171 vdd.t385 574.104
R608 vdd.t26 vdd.t47 574.104
R609 vdd.t450 vdd.t192 574.104
R610 vdd.t109 vdd.t368 574.104
R611 vdd.t179 vdd.t264 574.104
R612 vdd.t339 vdd.t322 574.104
R613 vdd.t130 vdd.t140 574.104
R614 vdd.t126 vdd.t481 574.104
R615 vdd.t404 vdd.t514 574.104
R616 vdd.t169 vdd.t29 574.104
R617 vdd.t166 vdd.t160 574.104
R618 vdd.t370 vdd.t270 574.104
R619 vdd.t444 vdd.t65 574.104
R620 vdd.t149 vdd.t382 574.104
R621 vdd.t86 vdd.t40 574.104
R622 vdd.t155 vdd.t112 574.104
R623 vdd.t293 vdd.t53 574.104
R624 vdd.n98 vdd.t502 569.302
R625 vdd.n61 vdd.t289 564.744
R626 vdd.n54 vdd.t90 564.744
R627 vdd.n47 vdd.t267 564.744
R628 vdd.n40 vdd.t50 564.744
R629 vdd.n33 vdd.t11 564.744
R630 vdd.n26 vdd.t36 564.744
R631 vdd.n19 vdd.t96 564.744
R632 vdd.n12 vdd.t242 564.744
R633 vdd.n5 vdd.t469 564.744
R634 vdd.n62 vdd.n61 474.26
R635 vdd.n55 vdd.n54 474.26
R636 vdd.n48 vdd.n47 474.26
R637 vdd.n41 vdd.n40 474.26
R638 vdd.n34 vdd.n33 474.26
R639 vdd.n27 vdd.n26 474.26
R640 vdd.n20 vdd.n19 474.26
R641 vdd.n13 vdd.n12 474.26
R642 vdd.n6 vdd.n5 474.26
R643 vdd.n65 vdd.t375 471.139
R644 vdd.n58 vdd.t103 471.139
R645 vdd.n51 vdd.t13 471.139
R646 vdd.n44 vdd.t363 471.139
R647 vdd.n37 vdd.t319 471.139
R648 vdd.n30 vdd.t457 471.139
R649 vdd.n23 vdd.t533 471.139
R650 vdd.n16 vdd.t411 471.139
R651 vdd.n9 vdd.t440 471.139
R652 vdd.n2 vdd.t114 471.139
R653 vdd vdd.t137 410.296
R654 vdd vdd.t473 410.296
R655 vdd vdd.t121 410.296
R656 vdd vdd.t492 410.296
R657 vdd vdd.t145 410.296
R658 vdd vdd.t425 410.296
R659 vdd vdd.t461 410.296
R660 vdd vdd.t436 410.296
R661 vdd vdd.t94 410.296
R662 vdd vdd.t185 410.296
R663 vdd.t393 vdd.t521 405.616
R664 vdd.t500 vdd.t274 405.616
R665 vdd.t195 vdd.t31 405.616
R666 vdd.t385 vdd.t279 405.616
R667 vdd.t47 vdd.t527 405.616
R668 vdd.t192 vdd.t281 405.616
R669 vdd.t368 vdd.t223 405.616
R670 vdd.t264 vdd.t272 405.616
R671 vdd.t322 vdd.t33 405.616
R672 vdd.t140 vdd.t335 405.616
R673 vdd.t481 vdd.t525 405.616
R674 vdd.t514 vdd.t304 405.616
R675 vdd.t29 vdd.t519 405.616
R676 vdd.t160 vdd.t306 405.616
R677 vdd.t270 vdd.t254 405.616
R678 vdd.t65 vdd.t285 405.616
R679 vdd.t382 vdd.t256 405.616
R680 vdd.t40 vdd.t283 405.616
R681 vdd.t112 vdd.t523 405.616
R682 vdd.t53 vdd.t287 405.616
R683 vdd vdd.t510 390.017
R684 vdd vdd.t512 390.017
R685 vdd vdd.t55 390.017
R686 vdd vdd.t2 390.017
R687 vdd vdd.t38 390.017
R688 vdd vdd.t231 390.017
R689 vdd vdd.t0 390.017
R690 vdd vdd.t189 390.017
R691 vdd vdd.t233 390.017
R692 vdd vdd.t508 390.017
R693 vdd.t128 vdd.t57 374.416
R694 vdd.t438 vdd.t415 374.416
R695 vdd.t262 vdd.t315 374.416
R696 vdd.t517 vdd.t427 374.416
R697 vdd.t489 vdd.t139 374.416
R698 vdd.t379 vdd.t44 374.416
R699 vdd.t157 vdd.t35 374.416
R700 vdd.t413 vdd.t316 374.416
R701 vdd.t448 vdd.t153 374.416
R702 vdd.t175 vdd.t100 374.416
R703 vdd.t98 vdd.t168 374.416
R704 vdd.t475 vdd.t147 374.416
R705 vdd.t119 vdd.t374 374.416
R706 vdd.t181 vdd.t387 374.416
R707 vdd.t372 vdd.t125 374.416
R708 vdd.t58 vdd.t191 374.416
R709 vdd.t151 vdd.t148 374.416
R710 vdd.t428 vdd.t454 374.416
R711 vdd.t6 vdd.t134 374.416
R712 vdd.t4 vdd.t23 374.416
R713 vdd.t510 vdd.t430 318.253
R714 vdd.t135 vdd.t128 318.253
R715 vdd.t57 vdd.t392 318.253
R716 vdd.t377 vdd.t438 318.253
R717 vdd.t415 vdd.t499 318.253
R718 vdd.t512 vdd.t418 318.253
R719 vdd.t471 vdd.t262 318.253
R720 vdd.t315 vdd.t197 318.253
R721 vdd.t101 vdd.t517 318.253
R722 vdd.t427 vdd.t384 318.253
R723 vdd.t55 vdd.t173 318.253
R724 vdd.t123 vdd.t489 318.253
R725 vdd.t139 vdd.t49 318.253
R726 vdd.t15 vdd.t379 318.253
R727 vdd.t44 vdd.t194 318.253
R728 vdd.t2 vdd.t452 318.253
R729 vdd.t494 vdd.t157 318.253
R730 vdd.t35 vdd.t367 318.253
R731 vdd.t365 vdd.t413 318.253
R732 vdd.t316 vdd.t266 318.253
R733 vdd.t38 vdd.t177 318.253
R734 vdd.t143 vdd.t448 318.253
R735 vdd.t153 vdd.t321 318.253
R736 vdd.t317 vdd.t175 318.253
R737 vdd.t100 vdd.t142 318.253
R738 vdd.t231 vdd.t132 318.253
R739 vdd.t423 vdd.t98 318.253
R740 vdd.t168 vdd.t483 318.253
R741 vdd.t455 vdd.t475 318.253
R742 vdd.t147 vdd.t516 318.253
R743 vdd.t0 vdd.t406 318.253
R744 vdd.t459 vdd.t119 318.253
R745 vdd.t374 vdd.t28 318.253
R746 vdd.t535 vdd.t181 318.253
R747 vdd.t387 vdd.t159 318.253
R748 vdd.t189 vdd.t164 318.253
R749 vdd.t434 vdd.t372 318.253
R750 vdd.t125 vdd.t269 318.253
R751 vdd.t409 vdd.t58 318.253
R752 vdd.t191 vdd.t67 318.253
R753 vdd.t233 vdd.t446 318.253
R754 vdd.t92 vdd.t151 318.253
R755 vdd.t148 vdd.t381 318.253
R756 vdd.t442 vdd.t428 318.253
R757 vdd.t454 vdd.t42 318.253
R758 vdd.t508 vdd.t88 318.253
R759 vdd.t183 vdd.t6 318.253
R760 vdd.t134 vdd.t111 318.253
R761 vdd.t116 vdd.t4 318.253
R762 vdd.t23 vdd.t52 318.253
R763 vdd.n237 vdd 293.171
R764 vdd vdd.n65 288.613
R765 vdd vdd.n62 288.613
R766 vdd vdd.n58 288.613
R767 vdd vdd.n55 288.613
R768 vdd vdd.n51 288.613
R769 vdd vdd.n48 288.613
R770 vdd vdd.n44 288.613
R771 vdd vdd.n41 288.613
R772 vdd vdd.n37 288.613
R773 vdd vdd.n34 288.613
R774 vdd vdd.n30 288.613
R775 vdd vdd.n27 288.613
R776 vdd vdd.n23 288.613
R777 vdd vdd.n20 288.613
R778 vdd vdd.n16 288.613
R779 vdd vdd.n13 288.613
R780 vdd vdd.n9 288.613
R781 vdd vdd.n6 288.613
R782 vdd vdd.n2 288.613
R783 vdd.n70 vdd.t390 242.278
R784 vdd.n73 vdd.t487 242.278
R785 vdd.n76 vdd.t188 242.278
R786 vdd.n79 vdd.t201 242.278
R787 vdd.n82 vdd.t538 242.278
R788 vdd.n85 vdd.t216 242.278
R789 vdd.n88 vdd.t85 242.278
R790 vdd.n91 vdd.t485 242.278
R791 vdd.n94 vdd.t432 242.278
R792 vdd.n97 vdd.t328 242.278
R793 vdd.t392 vdd.t397 230.889
R794 vdd.t499 vdd.t416 230.889
R795 vdd.t197 vdd.t105 230.889
R796 vdd.t384 vdd.t171 230.889
R797 vdd.t49 vdd.t26 230.889
R798 vdd.t194 vdd.t450 230.889
R799 vdd.t367 vdd.t109 230.889
R800 vdd.t266 vdd.t179 230.889
R801 vdd.t321 vdd.t339 230.889
R802 vdd.t142 vdd.t130 230.889
R803 vdd.t483 vdd.t126 230.889
R804 vdd.t516 vdd.t404 230.889
R805 vdd.t28 vdd.t169 230.889
R806 vdd.t159 vdd.t166 230.889
R807 vdd.t269 vdd.t370 230.889
R808 vdd.t67 vdd.t444 230.889
R809 vdd.t381 vdd.t149 230.889
R810 vdd.t42 vdd.t86 230.889
R811 vdd.t111 vdd.t155 230.889
R812 vdd.t52 vdd.t293 230.889
R813 vdd.t229 vdd 195.008
R814 vdd.t395 vdd 195.008
R815 vdd.t107 vdd 195.008
R816 vdd.t496 vdd 195.008
R817 vdd.t21 vdd 195.008
R818 vdd.t63 vdd 195.008
R819 vdd.t45 vdd 195.008
R820 vdd.t240 vdd 195.008
R821 vdd.t399 vdd 195.008
R822 vdd.t24 vdd 195.008
R823 vdd.t502 vdd 195.008
R824 vdd.t521 vdd 195.008
R825 vdd.t274 vdd 195.008
R826 vdd.t289 vdd 195.008
R827 vdd.t31 vdd 195.008
R828 vdd.t279 vdd 195.008
R829 vdd.t90 vdd 195.008
R830 vdd.t527 vdd 195.008
R831 vdd.t281 vdd 195.008
R832 vdd.t267 vdd 195.008
R833 vdd.t223 vdd 195.008
R834 vdd.t272 vdd 195.008
R835 vdd.t50 vdd 195.008
R836 vdd.t33 vdd 195.008
R837 vdd.t335 vdd 195.008
R838 vdd.t11 vdd 195.008
R839 vdd.t525 vdd 195.008
R840 vdd.t304 vdd 195.008
R841 vdd.t36 vdd 195.008
R842 vdd.t519 vdd 195.008
R843 vdd.t306 vdd 195.008
R844 vdd.t96 vdd 195.008
R845 vdd.t254 vdd 195.008
R846 vdd.t285 vdd 195.008
R847 vdd.t242 vdd 195.008
R848 vdd.t256 vdd 195.008
R849 vdd.t283 vdd 195.008
R850 vdd.t469 vdd 195.008
R851 vdd.t523 vdd 195.008
R852 vdd.t287 vdd 195.008
R853 vdd.t430 vdd 165.368
R854 vdd.t418 vdd 165.368
R855 vdd.t173 vdd 165.368
R856 vdd.t452 vdd 165.368
R857 vdd.t177 vdd 165.368
R858 vdd.t132 vdd 165.368
R859 vdd.t406 vdd 165.368
R860 vdd.t164 vdd 165.368
R861 vdd.t446 vdd 165.368
R862 vdd.t88 vdd 165.368
R863 vdd.t390 vdd.t246 148.7
R864 vdd.t246 vdd.t244 148.7
R865 vdd.t244 vdd.t389 148.7
R866 vdd.t389 vdd.t331 148.7
R867 vdd.t331 vdd.t402 148.7
R868 vdd.t402 vdd.t203 148.7
R869 vdd.t203 vdd.t504 148.7
R870 vdd.t504 vdd.t313 148.7
R871 vdd.t313 vdd.t245 148.7
R872 vdd.t245 vdd.t391 148.7
R873 vdd.t391 vdd.t312 148.7
R874 vdd.t312 vdd.t330 148.7
R875 vdd.t330 vdd.t401 148.7
R876 vdd.t401 vdd.t506 148.7
R877 vdd.t506 vdd.t314 148.7
R878 vdd.t314 vdd.t204 148.7
R879 vdd.t204 vdd.t505 148.7
R880 vdd.t487 vdd.t309 148.7
R881 vdd.t309 vdd.t354 148.7
R882 vdd.t354 vdd.t347 148.7
R883 vdd.t347 vdd.t356 148.7
R884 vdd.t356 vdd.t338 148.7
R885 vdd.t338 vdd.t301 148.7
R886 vdd.t301 vdd.t488 148.7
R887 vdd.t488 vdd.t261 148.7
R888 vdd.t261 vdd.t299 148.7
R889 vdd.t299 vdd.t348 148.7
R890 vdd.t348 vdd.t357 148.7
R891 vdd.t357 vdd.t355 148.7
R892 vdd.t355 vdd.t337 148.7
R893 vdd.t337 vdd.t300 148.7
R894 vdd.t300 vdd.t341 148.7
R895 vdd.t341 vdd.t308 148.7
R896 vdd.t308 vdd.t349 148.7
R897 vdd.t188 vdd.t303 148.7
R898 vdd.t303 vdd.t353 148.7
R899 vdd.t353 vdd.t403 148.7
R900 vdd.t403 vdd.t278 148.7
R901 vdd.t278 vdd.t239 148.7
R902 vdd.t239 vdd.t163 148.7
R903 vdd.t163 vdd.t162 148.7
R904 vdd.t162 vdd.t238 148.7
R905 vdd.t238 vdd.t292 148.7
R906 vdd.t292 vdd.t334 148.7
R907 vdd.t334 vdd.t187 148.7
R908 vdd.t187 vdd.t507 148.7
R909 vdd.t507 vdd.t333 148.7
R910 vdd.t333 vdd.t491 148.7
R911 vdd.t491 vdd.t209 148.7
R912 vdd.t209 vdd.t302 148.7
R913 vdd.t302 vdd.t352 148.7
R914 vdd.t201 vdd.t199 148.7
R915 vdd.t199 vdd.t250 148.7
R916 vdd.t250 vdd.t200 148.7
R917 vdd.t200 vdd.t198 148.7
R918 vdd.t198 vdd.t247 148.7
R919 vdd.t247 vdd.t212 148.7
R920 vdd.t212 vdd.t360 148.7
R921 vdd.t360 vdd.t214 148.7
R922 vdd.t214 vdd.t154 148.7
R923 vdd.t154 vdd.t202 148.7
R924 vdd.t202 vdd.t362 148.7
R925 vdd.t362 vdd.t249 148.7
R926 vdd.t249 vdd.t205 148.7
R927 vdd.t205 vdd.t361 148.7
R928 vdd.t361 vdd.t248 148.7
R929 vdd.t248 vdd.t213 148.7
R930 vdd.t213 vdd.t206 148.7
R931 vdd.t538 vdd.t9 148.7
R932 vdd.t9 vdd.t226 148.7
R933 vdd.t226 vdd.t537 148.7
R934 vdd.t537 vdd.t8 148.7
R935 vdd.t8 vdd.t235 148.7
R936 vdd.t235 vdd.t228 148.7
R937 vdd.t228 vdd.t62 148.7
R938 vdd.t62 vdd.t60 148.7
R939 vdd.t60 vdd.t227 148.7
R940 vdd.t227 vdd.t539 148.7
R941 vdd.t539 vdd.t10 148.7
R942 vdd.t10 vdd.t236 148.7
R943 vdd.t236 vdd.t332 148.7
R944 vdd.t332 vdd.t277 148.7
R945 vdd.t277 vdd.t61 148.7
R946 vdd.t61 vdd.t225 148.7
R947 vdd.t225 vdd.t276 148.7
R948 vdd.t216 vdd.t251 148.7
R949 vdd.t251 vdd.t220 148.7
R950 vdd.t220 vdd.t388 148.7
R951 vdd.t388 vdd.t207 148.7
R952 vdd.t207 vdd.t219 148.7
R953 vdd.t219 vdd.t208 148.7
R954 vdd.t208 vdd.t217 148.7
R955 vdd.t217 vdd.t253 148.7
R956 vdd.t253 vdd.t222 148.7
R957 vdd.t222 vdd.t258 148.7
R958 vdd.t258 vdd.t252 148.7
R959 vdd.t252 vdd.t221 148.7
R960 vdd.t221 vdd.t237 148.7
R961 vdd.t237 vdd.t260 148.7
R962 vdd.t260 vdd.t215 148.7
R963 vdd.t215 vdd.t218 148.7
R964 vdd.t218 vdd.t259 148.7
R965 vdd.t85 vdd.t69 148.7
R966 vdd.t69 vdd.t78 148.7
R967 vdd.t78 vdd.t75 148.7
R968 vdd.t75 vdd.t82 148.7
R969 vdd.t82 vdd.t72 148.7
R970 vdd.t72 vdd.t76 148.7
R971 vdd.t76 vdd.t83 148.7
R972 vdd.t83 vdd.t68 148.7
R973 vdd.t68 vdd.t70 148.7
R974 vdd.t70 vdd.t79 148.7
R975 vdd.t79 vdd.t80 148.7
R976 vdd.t80 vdd.t71 148.7
R977 vdd.t71 vdd.t74 148.7
R978 vdd.t74 vdd.t81 148.7
R979 vdd.t81 vdd.t73 148.7
R980 vdd.t73 vdd.t77 148.7
R981 vdd.t77 vdd.t84 148.7
R982 vdd.t485 vdd.t18 148.7
R983 vdd.t18 vdd.t17 148.7
R984 vdd.t17 vdd.t532 148.7
R985 vdd.t532 vdd.t484 148.7
R986 vdd.t484 vdd.t468 148.7
R987 vdd.t468 vdd.t463 148.7
R988 vdd.t463 vdd.t19 148.7
R989 vdd.t19 vdd.t467 148.7
R990 vdd.t467 vdd.t20 148.7
R991 vdd.t20 vdd.t486 148.7
R992 vdd.t486 vdd.t531 148.7
R993 vdd.t531 vdd.t478 148.7
R994 vdd.t478 vdd.t465 148.7
R995 vdd.t465 vdd.t43 148.7
R996 vdd.t43 vdd.t477 148.7
R997 vdd.t477 vdd.t464 148.7
R998 vdd.t464 vdd.t466 148.7
R999 vdd.t432 vdd.t118 148.7
R1000 vdd.t118 vdd.t291 148.7
R1001 vdd.t291 vdd.t480 148.7
R1002 vdd.t480 vdd.t359 148.7
R1003 vdd.t359 vdd.t530 148.7
R1004 vdd.t530 vdd.t311 148.7
R1005 vdd.t311 vdd.t342 148.7
R1006 vdd.t342 vdd.t421 148.7
R1007 vdd.t421 vdd.t310 148.7
R1008 vdd.t310 vdd.t433 148.7
R1009 vdd.t433 vdd.t479 148.7
R1010 vdd.t479 vdd.t358 148.7
R1011 vdd.t358 vdd.t529 148.7
R1012 vdd.t529 vdd.t351 148.7
R1013 vdd.t351 vdd.t422 148.7
R1014 vdd.t422 vdd.t420 148.7
R1015 vdd.t420 vdd.t350 148.7
R1016 vdd.t328 vdd.t295 148.7
R1017 vdd.t295 vdd.t498 148.7
R1018 vdd.t498 vdd.t324 148.7
R1019 vdd.t324 vdd.t345 148.7
R1020 vdd.t345 vdd.t210 148.7
R1021 vdd.t210 vdd.t325 148.7
R1022 vdd.t325 vdd.t211 148.7
R1023 vdd.t211 vdd.t297 148.7
R1024 vdd.t297 vdd.t326 148.7
R1025 vdd.t326 vdd.t343 148.7
R1026 vdd.t343 vdd.t346 148.7
R1027 vdd.t346 vdd.t329 148.7
R1028 vdd.t329 vdd.t296 148.7
R1029 vdd.t296 vdd.t344 148.7
R1030 vdd.t344 vdd.t298 148.7
R1031 vdd.t298 vdd.t327 148.7
R1032 vdd.t327 vdd.t408 148.7
R1033 vdd.n226 vdd.t509 15.5636
R1034 vdd.n212 vdd.t234 15.5636
R1035 vdd.n198 vdd.t190 15.5636
R1036 vdd.n184 vdd.t1 15.5636
R1037 vdd.n170 vdd.t232 15.5636
R1038 vdd.n156 vdd.t39 15.5636
R1039 vdd.n142 vdd.t3 15.5636
R1040 vdd.n128 vdd.t56 15.5636
R1041 vdd.n114 vdd.t513 15.5636
R1042 vdd.n100 vdd.t511 15.5636
R1043 vdd.n235 vdd.t294 4.77854
R1044 vdd.n230 vdd.t156 4.77854
R1045 vdd.n221 vdd.t87 4.77854
R1046 vdd.n216 vdd.t150 4.77854
R1047 vdd.n207 vdd.t445 4.77854
R1048 vdd.n202 vdd.t371 4.77854
R1049 vdd.n193 vdd.t167 4.77854
R1050 vdd.n188 vdd.t170 4.77854
R1051 vdd.n179 vdd.t405 4.77854
R1052 vdd.n174 vdd.t127 4.77854
R1053 vdd.n165 vdd.t131 4.77854
R1054 vdd.n160 vdd.t340 4.77854
R1055 vdd.n151 vdd.t180 4.77854
R1056 vdd.n146 vdd.t110 4.77854
R1057 vdd.n137 vdd.t451 4.77854
R1058 vdd.n132 vdd.t27 4.77854
R1059 vdd.n123 vdd.t172 4.77854
R1060 vdd.n118 vdd.t106 4.77854
R1061 vdd.n109 vdd.t417 4.77854
R1062 vdd.n104 vdd.t398 4.77854
R1063 vdd.n98 vdd.n97 4.69929
R1064 vdd.n232 vdd.n2 4.55932
R1065 vdd.n224 vdd.n5 4.55932
R1066 vdd.n223 vdd.n6 4.55932
R1067 vdd.n218 vdd.n9 4.55932
R1068 vdd.n210 vdd.n12 4.55932
R1069 vdd.n209 vdd.n13 4.55932
R1070 vdd.n204 vdd.n16 4.55932
R1071 vdd.n196 vdd.n19 4.55932
R1072 vdd.n195 vdd.n20 4.55932
R1073 vdd.n190 vdd.n23 4.55932
R1074 vdd.n182 vdd.n26 4.55932
R1075 vdd.n181 vdd.n27 4.55932
R1076 vdd.n176 vdd.n30 4.55932
R1077 vdd.n168 vdd.n33 4.55932
R1078 vdd.n167 vdd.n34 4.55932
R1079 vdd.n162 vdd.n37 4.55932
R1080 vdd.n154 vdd.n40 4.55932
R1081 vdd.n153 vdd.n41 4.55932
R1082 vdd.n148 vdd.n44 4.55932
R1083 vdd.n140 vdd.n47 4.55932
R1084 vdd.n139 vdd.n48 4.55932
R1085 vdd.n134 vdd.n51 4.55932
R1086 vdd.n126 vdd.n54 4.55932
R1087 vdd.n125 vdd.n55 4.55932
R1088 vdd.n120 vdd.n58 4.55932
R1089 vdd.n112 vdd.n61 4.55932
R1090 vdd.n111 vdd.n62 4.55932
R1091 vdd.n106 vdd.n65 4.55932
R1092 vdd.n233 vdd.t115 3.95308
R1093 vdd.n228 vdd.t186 3.95308
R1094 vdd.n219 vdd.t441 3.95308
R1095 vdd.n214 vdd.t95 3.95308
R1096 vdd.n205 vdd.t412 3.95308
R1097 vdd.n200 vdd.t437 3.95308
R1098 vdd.n191 vdd.t534 3.95308
R1099 vdd.n186 vdd.t462 3.95308
R1100 vdd.n177 vdd.t458 3.95308
R1101 vdd.n172 vdd.t426 3.95308
R1102 vdd.n163 vdd.t320 3.95308
R1103 vdd.n158 vdd.t146 3.95308
R1104 vdd.n149 vdd.t364 3.95308
R1105 vdd.n144 vdd.t493 3.95308
R1106 vdd.n135 vdd.t14 3.95308
R1107 vdd.n130 vdd.t122 3.95308
R1108 vdd.n121 vdd.t104 3.95308
R1109 vdd.n116 vdd.t474 3.95308
R1110 vdd.n107 vdd.t376 3.95308
R1111 vdd.n102 vdd.t138 3.95308
R1112 vdd.n227 vdd.t89 3.90058
R1113 vdd.n213 vdd.t447 3.90058
R1114 vdd.n199 vdd.t165 3.90058
R1115 vdd.n185 vdd.t407 3.90058
R1116 vdd.n171 vdd.t133 3.90058
R1117 vdd.n157 vdd.t178 3.90058
R1118 vdd.n143 vdd.t453 3.90058
R1119 vdd.n129 vdd.t174 3.90058
R1120 vdd.n115 vdd.t419 3.90058
R1121 vdd.n101 vdd.t431 3.90058
R1122 vdd.n69 vdd.t230 3.84351
R1123 vdd.n72 vdd.t396 3.84351
R1124 vdd.n75 vdd.t108 3.84351
R1125 vdd.n78 vdd.t497 3.84351
R1126 vdd.n81 vdd.t22 3.84351
R1127 vdd.n84 vdd.t64 3.84351
R1128 vdd.n87 vdd.t46 3.84351
R1129 vdd.n90 vdd.t241 3.84351
R1130 vdd.n93 vdd.t400 3.84351
R1131 vdd.n96 vdd.t25 3.84351
R1132 vdd.n225 vdd.t470 3.84351
R1133 vdd.n211 vdd.t243 3.84351
R1134 vdd.n197 vdd.t97 3.84351
R1135 vdd.n183 vdd.t37 3.84351
R1136 vdd.n169 vdd.t12 3.84351
R1137 vdd.n155 vdd.t51 3.84351
R1138 vdd.n141 vdd.t268 3.84351
R1139 vdd.n127 vdd.t91 3.84351
R1140 vdd.n113 vdd.t290 3.84351
R1141 vdd.n99 vdd.t503 3.84351
R1142 vdd.n0 vdd.t54 3.7805
R1143 vdd.n3 vdd.t113 3.7805
R1144 vdd.n7 vdd.t41 3.7805
R1145 vdd.n10 vdd.t383 3.7805
R1146 vdd.n14 vdd.t66 3.7805
R1147 vdd.n17 vdd.t271 3.7805
R1148 vdd.n21 vdd.t161 3.7805
R1149 vdd.n24 vdd.t30 3.7805
R1150 vdd.n28 vdd.t515 3.7805
R1151 vdd.n31 vdd.t482 3.7805
R1152 vdd.n35 vdd.t141 3.7805
R1153 vdd.n38 vdd.t323 3.7805
R1154 vdd.n42 vdd.t265 3.7805
R1155 vdd.n45 vdd.t369 3.7805
R1156 vdd.n49 vdd.t193 3.7805
R1157 vdd.n52 vdd.t48 3.7805
R1158 vdd.n56 vdd.t386 3.7805
R1159 vdd.n59 vdd.t196 3.7805
R1160 vdd.n63 vdd.t501 3.7805
R1161 vdd.n66 vdd.t394 3.7805
R1162 vdd.n73 vdd.n72 3.0298
R1163 vdd.n76 vdd.n75 3.0298
R1164 vdd.n79 vdd.n78 3.0298
R1165 vdd.n82 vdd.n81 3.0298
R1166 vdd.n85 vdd.n84 3.0298
R1167 vdd.n88 vdd.n87 3.0298
R1168 vdd.n91 vdd.n90 3.0298
R1169 vdd.n94 vdd.n93 3.0298
R1170 vdd.n97 vdd.n96 3.0298
R1171 vdd.n236 vdd.n0 2.95854
R1172 vdd.n234 vdd.n1 2.95854
R1173 vdd.n231 vdd.n3 2.95854
R1174 vdd.n229 vdd.n4 2.95854
R1175 vdd.n222 vdd.n7 2.95854
R1176 vdd.n220 vdd.n8 2.95854
R1177 vdd.n217 vdd.n10 2.95854
R1178 vdd.n215 vdd.n11 2.95854
R1179 vdd.n208 vdd.n14 2.95854
R1180 vdd.n206 vdd.n15 2.95854
R1181 vdd.n203 vdd.n17 2.95854
R1182 vdd.n201 vdd.n18 2.95854
R1183 vdd.n194 vdd.n21 2.95854
R1184 vdd.n192 vdd.n22 2.95854
R1185 vdd.n189 vdd.n24 2.95854
R1186 vdd.n187 vdd.n25 2.95854
R1187 vdd.n180 vdd.n28 2.95854
R1188 vdd.n178 vdd.n29 2.95854
R1189 vdd.n175 vdd.n31 2.95854
R1190 vdd.n173 vdd.n32 2.95854
R1191 vdd.n166 vdd.n35 2.95854
R1192 vdd.n164 vdd.n36 2.95854
R1193 vdd.n161 vdd.n38 2.95854
R1194 vdd.n159 vdd.n39 2.95854
R1195 vdd.n152 vdd.n42 2.95854
R1196 vdd.n150 vdd.n43 2.95854
R1197 vdd.n147 vdd.n45 2.95854
R1198 vdd.n145 vdd.n46 2.95854
R1199 vdd.n138 vdd.n49 2.95854
R1200 vdd.n136 vdd.n50 2.95854
R1201 vdd.n133 vdd.n52 2.95854
R1202 vdd.n131 vdd.n53 2.95854
R1203 vdd.n124 vdd.n56 2.95854
R1204 vdd.n122 vdd.n57 2.95854
R1205 vdd.n119 vdd.n59 2.95854
R1206 vdd.n117 vdd.n60 2.95854
R1207 vdd.n110 vdd.n63 2.95854
R1208 vdd.n108 vdd.n64 2.95854
R1209 vdd.n105 vdd.n66 2.95854
R1210 vdd.n103 vdd.n67 2.95854
R1211 vdd.n70 vdd.n69 2.84768
R1212 vdd.n0 vdd.t288 1.53332
R1213 vdd.n3 vdd.t524 1.53332
R1214 vdd.n7 vdd.t284 1.53332
R1215 vdd.n10 vdd.t257 1.53332
R1216 vdd.n14 vdd.t286 1.53332
R1217 vdd.n17 vdd.t255 1.53332
R1218 vdd.n21 vdd.t307 1.53332
R1219 vdd.n24 vdd.t520 1.53332
R1220 vdd.n28 vdd.t305 1.53332
R1221 vdd.n31 vdd.t526 1.53332
R1222 vdd.n35 vdd.t336 1.53332
R1223 vdd.n38 vdd.t34 1.53332
R1224 vdd.n42 vdd.t273 1.53332
R1225 vdd.n45 vdd.t224 1.53332
R1226 vdd.n49 vdd.t282 1.53332
R1227 vdd.n52 vdd.t528 1.53332
R1228 vdd.n56 vdd.t280 1.53332
R1229 vdd.n59 vdd.t32 1.53332
R1230 vdd.n63 vdd.t275 1.53332
R1231 vdd.n66 vdd.t522 1.53332
R1232 vdd.n1 vdd.t117 1.31934
R1233 vdd.n1 vdd.t5 1.31934
R1234 vdd.n4 vdd.t184 1.31934
R1235 vdd.n4 vdd.t7 1.31934
R1236 vdd.n8 vdd.t443 1.31934
R1237 vdd.n8 vdd.t429 1.31934
R1238 vdd.n11 vdd.t93 1.31934
R1239 vdd.n11 vdd.t152 1.31934
R1240 vdd.n15 vdd.t410 1.31934
R1241 vdd.n15 vdd.t59 1.31934
R1242 vdd.n18 vdd.t435 1.31934
R1243 vdd.n18 vdd.t373 1.31934
R1244 vdd.n22 vdd.t536 1.31934
R1245 vdd.n22 vdd.t182 1.31934
R1246 vdd.n25 vdd.t460 1.31934
R1247 vdd.n25 vdd.t120 1.31934
R1248 vdd.n29 vdd.t456 1.31934
R1249 vdd.n29 vdd.t476 1.31934
R1250 vdd.n32 vdd.t424 1.31934
R1251 vdd.n32 vdd.t99 1.31934
R1252 vdd.n36 vdd.t318 1.31934
R1253 vdd.n36 vdd.t176 1.31934
R1254 vdd.n39 vdd.t144 1.31934
R1255 vdd.n39 vdd.t449 1.31934
R1256 vdd.n43 vdd.t366 1.31934
R1257 vdd.n43 vdd.t414 1.31934
R1258 vdd.n46 vdd.t495 1.31934
R1259 vdd.n46 vdd.t158 1.31934
R1260 vdd.n50 vdd.t16 1.31934
R1261 vdd.n50 vdd.t380 1.31934
R1262 vdd.n53 vdd.t124 1.31934
R1263 vdd.n53 vdd.t490 1.31934
R1264 vdd.n57 vdd.t102 1.31934
R1265 vdd.n57 vdd.t518 1.31934
R1266 vdd.n60 vdd.t472 1.31934
R1267 vdd.n60 vdd.t263 1.31934
R1268 vdd.n64 vdd.t378 1.31934
R1269 vdd.n64 vdd.t439 1.31934
R1270 vdd.n67 vdd.t136 1.31934
R1271 vdd.n67 vdd.t129 1.31934
R1272 vdd vdd.n70 0.614627
R1273 vdd vdd.n73 0.557603
R1274 vdd vdd.n76 0.557603
R1275 vdd vdd.n79 0.557603
R1276 vdd vdd.n82 0.557603
R1277 vdd vdd.n85 0.557603
R1278 vdd vdd.n88 0.557603
R1279 vdd vdd.n91 0.557603
R1280 vdd vdd.n94 0.557603
R1281 vdd.n104 vdd.n103 0.3985
R1282 vdd.n109 vdd.n108 0.3985
R1283 vdd.n118 vdd.n117 0.3985
R1284 vdd.n123 vdd.n122 0.3985
R1285 vdd.n132 vdd.n131 0.3985
R1286 vdd.n137 vdd.n136 0.3985
R1287 vdd.n146 vdd.n145 0.3985
R1288 vdd.n151 vdd.n150 0.3985
R1289 vdd.n160 vdd.n159 0.3985
R1290 vdd.n165 vdd.n164 0.3985
R1291 vdd.n174 vdd.n173 0.3985
R1292 vdd.n179 vdd.n178 0.3985
R1293 vdd.n188 vdd.n187 0.3985
R1294 vdd.n193 vdd.n192 0.3985
R1295 vdd.n202 vdd.n201 0.3985
R1296 vdd.n207 vdd.n206 0.3985
R1297 vdd.n216 vdd.n215 0.3985
R1298 vdd.n221 vdd.n220 0.3985
R1299 vdd.n230 vdd.n229 0.3985
R1300 vdd.n235 vdd.n234 0.3985
R1301 vdd.n103 vdd.n102 0.3165
R1302 vdd.n108 vdd.n107 0.3165
R1303 vdd.n117 vdd.n116 0.3165
R1304 vdd.n122 vdd.n121 0.3165
R1305 vdd.n131 vdd.n130 0.3165
R1306 vdd.n136 vdd.n135 0.3165
R1307 vdd.n145 vdd.n144 0.3165
R1308 vdd.n150 vdd.n149 0.3165
R1309 vdd.n159 vdd.n158 0.3165
R1310 vdd.n164 vdd.n163 0.3165
R1311 vdd.n173 vdd.n172 0.3165
R1312 vdd.n178 vdd.n177 0.3165
R1313 vdd.n187 vdd.n186 0.3165
R1314 vdd.n192 vdd.n191 0.3165
R1315 vdd.n201 vdd.n200 0.3165
R1316 vdd.n206 vdd.n205 0.3165
R1317 vdd.n215 vdd.n214 0.3165
R1318 vdd.n220 vdd.n219 0.3165
R1319 vdd.n229 vdd.n228 0.3165
R1320 vdd.n234 vdd.n233 0.3165
R1321 vdd.n99 vdd.n98 0.2305
R1322 vdd.n113 vdd.n112 0.2305
R1323 vdd.n127 vdd.n126 0.2305
R1324 vdd.n141 vdd.n140 0.2305
R1325 vdd.n155 vdd.n154 0.2305
R1326 vdd.n169 vdd.n168 0.2305
R1327 vdd.n183 vdd.n182 0.2305
R1328 vdd.n197 vdd.n196 0.2305
R1329 vdd.n211 vdd.n210 0.2305
R1330 vdd.n225 vdd.n224 0.2305
R1331 vdd.n105 vdd.n104 0.2125
R1332 vdd.n110 vdd.n109 0.2125
R1333 vdd.n119 vdd.n118 0.2125
R1334 vdd.n124 vdd.n123 0.2125
R1335 vdd.n133 vdd.n132 0.2125
R1336 vdd.n138 vdd.n137 0.2125
R1337 vdd.n147 vdd.n146 0.2125
R1338 vdd.n152 vdd.n151 0.2125
R1339 vdd.n161 vdd.n160 0.2125
R1340 vdd.n166 vdd.n165 0.2125
R1341 vdd.n175 vdd.n174 0.2125
R1342 vdd.n180 vdd.n179 0.2125
R1343 vdd.n189 vdd.n188 0.2125
R1344 vdd.n194 vdd.n193 0.2125
R1345 vdd.n203 vdd.n202 0.2125
R1346 vdd.n208 vdd.n207 0.2125
R1347 vdd.n217 vdd.n216 0.2125
R1348 vdd.n222 vdd.n221 0.2125
R1349 vdd.n231 vdd.n230 0.2125
R1350 vdd.n236 vdd.n235 0.2125
R1351 vdd.n106 vdd.n105 0.2085
R1352 vdd.n120 vdd.n119 0.2085
R1353 vdd.n134 vdd.n133 0.2085
R1354 vdd.n148 vdd.n147 0.2085
R1355 vdd.n162 vdd.n161 0.2085
R1356 vdd.n176 vdd.n175 0.2085
R1357 vdd.n190 vdd.n189 0.2085
R1358 vdd.n204 vdd.n203 0.2085
R1359 vdd.n218 vdd.n217 0.2085
R1360 vdd.n232 vdd.n231 0.2085
R1361 vdd.n101 vdd.n100 0.2045
R1362 vdd.n115 vdd.n114 0.2045
R1363 vdd.n129 vdd.n128 0.2045
R1364 vdd.n143 vdd.n142 0.2045
R1365 vdd.n157 vdd.n156 0.2045
R1366 vdd.n171 vdd.n170 0.2045
R1367 vdd.n185 vdd.n184 0.2045
R1368 vdd.n199 vdd.n198 0.2045
R1369 vdd.n213 vdd.n212 0.2045
R1370 vdd.n227 vdd.n226 0.2045
R1371 vdd.n111 vdd 0.1415
R1372 vdd.n125 vdd 0.1415
R1373 vdd.n139 vdd 0.1415
R1374 vdd.n153 vdd 0.1415
R1375 vdd.n167 vdd 0.1415
R1376 vdd.n181 vdd 0.1415
R1377 vdd.n195 vdd 0.1415
R1378 vdd.n209 vdd 0.1415
R1379 vdd.n223 vdd 0.1415
R1380 vdd.n237 vdd 0.1415
R1381 vdd.n107 vdd.n106 0.0985
R1382 vdd.n121 vdd.n120 0.0985
R1383 vdd.n135 vdd.n134 0.0985
R1384 vdd.n149 vdd.n148 0.0985
R1385 vdd.n163 vdd.n162 0.0985
R1386 vdd.n177 vdd.n176 0.0985
R1387 vdd.n191 vdd.n190 0.0985
R1388 vdd.n205 vdd.n204 0.0985
R1389 vdd.n219 vdd.n218 0.0985
R1390 vdd.n233 vdd.n232 0.0985
R1391 vdd vdd.n71 0.0919062
R1392 vdd vdd.n74 0.0919062
R1393 vdd vdd.n77 0.0919062
R1394 vdd vdd.n80 0.0919062
R1395 vdd vdd.n83 0.0919062
R1396 vdd vdd.n86 0.0919062
R1397 vdd vdd.n89 0.0919062
R1398 vdd vdd.n92 0.0919062
R1399 vdd vdd.n95 0.0919062
R1400 vdd vdd.n68 0.0894058
R1401 vdd.n100 vdd.n99 0.086
R1402 vdd.n114 vdd.n113 0.086
R1403 vdd.n128 vdd.n127 0.086
R1404 vdd.n142 vdd.n141 0.086
R1405 vdd.n156 vdd.n155 0.086
R1406 vdd.n170 vdd.n169 0.086
R1407 vdd.n184 vdd.n183 0.086
R1408 vdd.n198 vdd.n197 0.086
R1409 vdd.n212 vdd.n211 0.086
R1410 vdd.n226 vdd.n225 0.086
R1411 vdd.n102 vdd.n101 0.083
R1412 vdd.n116 vdd.n115 0.083
R1413 vdd.n130 vdd.n129 0.083
R1414 vdd.n144 vdd.n143 0.083
R1415 vdd.n158 vdd.n157 0.083
R1416 vdd.n172 vdd.n171 0.083
R1417 vdd.n186 vdd.n185 0.083
R1418 vdd.n200 vdd.n199 0.083
R1419 vdd.n214 vdd.n213 0.083
R1420 vdd.n228 vdd.n227 0.083
R1421 vdd vdd.n111 0.0775
R1422 vdd vdd.n125 0.0775
R1423 vdd vdd.n139 0.0775
R1424 vdd vdd.n153 0.0775
R1425 vdd vdd.n167 0.0775
R1426 vdd vdd.n181 0.0775
R1427 vdd vdd.n195 0.0775
R1428 vdd vdd.n209 0.0775
R1429 vdd vdd.n223 0.0775
R1430 vdd vdd.n237 0.0775
R1431 vdd.n112 vdd 0.0755
R1432 vdd.n126 vdd 0.0755
R1433 vdd.n140 vdd 0.0755
R1434 vdd.n154 vdd 0.0755
R1435 vdd.n168 vdd 0.0755
R1436 vdd.n182 vdd 0.0755
R1437 vdd.n196 vdd 0.0755
R1438 vdd.n210 vdd 0.0755
R1439 vdd.n224 vdd 0.0755
R1440 vdd vdd.n110 0.0675
R1441 vdd vdd.n124 0.0675
R1442 vdd vdd.n138 0.0675
R1443 vdd vdd.n152 0.0675
R1444 vdd vdd.n166 0.0675
R1445 vdd vdd.n180 0.0675
R1446 vdd vdd.n194 0.0675
R1447 vdd vdd.n208 0.0675
R1448 vdd vdd.n222 0.0675
R1449 vdd vdd.n236 0.0675
R1450 vdd.n72 vdd 0.037625
R1451 vdd.n75 vdd 0.037625
R1452 vdd.n78 vdd 0.037625
R1453 vdd.n81 vdd 0.037625
R1454 vdd.n84 vdd 0.037625
R1455 vdd.n87 vdd 0.037625
R1456 vdd.n90 vdd 0.037625
R1457 vdd.n93 vdd 0.037625
R1458 vdd.n96 vdd 0.037625
R1459 vdd.n69 vdd 0.0366094
R1460 vdd.n71 vdd 0.001625
R1461 vdd.n74 vdd 0.001625
R1462 vdd.n77 vdd 0.001625
R1463 vdd.n80 vdd 0.001625
R1464 vdd.n83 vdd 0.001625
R1465 vdd.n86 vdd 0.001625
R1466 vdd.n89 vdd 0.001625
R1467 vdd.n92 vdd 0.001625
R1468 vdd.n95 vdd 0.001625
R1469 vdd.n68 vdd 0.00159422
R1470 BUS[2].n2 BUS[2].n0 15.3751
R1471 BUS[2].n9 BUS[2].n7 15.2168
R1472 BUS[2].n2 BUS[2].n1 15.0151
R1473 BUS[2].n4 BUS[2].n3 15.0151
R1474 BUS[2].n21 BUS[2].n20 14.8568
R1475 BUS[2].n19 BUS[2].n18 14.8568
R1476 BUS[2].n17 BUS[2].n16 14.8568
R1477 BUS[2].n15 BUS[2].n14 14.8568
R1478 BUS[2].n13 BUS[2].n12 14.8568
R1479 BUS[2].n11 BUS[2].n10 14.8568
R1480 BUS[2].n9 BUS[2].n8 14.8568
R1481 BUS[2].n6 BUS[2].n5 14.8568
R1482 BUS[2].n22 BUS[2] 0.921051
R1483 BUS[2].n6 BUS[2].n4 0.8825
R1484 BUS[2].n20 BUS[2].t2 0.4555
R1485 BUS[2].n20 BUS[2].t8 0.4555
R1486 BUS[2].n18 BUS[2].t13 0.4555
R1487 BUS[2].n18 BUS[2].t6 0.4555
R1488 BUS[2].n16 BUS[2].t10 0.4555
R1489 BUS[2].n16 BUS[2].t15 0.4555
R1490 BUS[2].n14 BUS[2].t0 0.4555
R1491 BUS[2].n14 BUS[2].t1 0.4555
R1492 BUS[2].n12 BUS[2].t3 0.4555
R1493 BUS[2].n12 BUS[2].t23 0.4555
R1494 BUS[2].n10 BUS[2].t14 0.4555
R1495 BUS[2].n10 BUS[2].t7 0.4555
R1496 BUS[2].n8 BUS[2].t12 0.4555
R1497 BUS[2].n8 BUS[2].t9 0.4555
R1498 BUS[2].n7 BUS[2].t22 0.4555
R1499 BUS[2].n7 BUS[2].t5 0.4555
R1500 BUS[2].n5 BUS[2].t4 0.4555
R1501 BUS[2].n5 BUS[2].t11 0.4555
R1502 BUS[2].n0 BUS[2].t17 0.41
R1503 BUS[2].n0 BUS[2].t20 0.41
R1504 BUS[2].n1 BUS[2].t19 0.41
R1505 BUS[2].n1 BUS[2].t16 0.41
R1506 BUS[2].n3 BUS[2].t21 0.41
R1507 BUS[2].n3 BUS[2].t18 0.41
R1508 BUS[2].n4 BUS[2].n2 0.3605
R1509 BUS[2].n11 BUS[2].n9 0.3605
R1510 BUS[2].n13 BUS[2].n11 0.3605
R1511 BUS[2].n15 BUS[2].n13 0.3605
R1512 BUS[2].n17 BUS[2].n15 0.3605
R1513 BUS[2].n19 BUS[2].n17 0.3605
R1514 BUS[2].n21 BUS[2].n19 0.3605
R1515 BUS[2].n22 BUS[2].n6 0.203
R1516 BUS[2] BUS[2].n22 0.0430197
R1517 BUS[2].n22 BUS[2].n21 0.015125
R1518 vss.n284 vss.n283 2.09667e+06
R1519 vss.t393 vss.n121 46438.4
R1520 vss.n118 vss.n117 42250
R1521 vss.n114 vss.n113 42250
R1522 vss.n110 vss.n109 42250
R1523 vss.n106 vss.n105 42250
R1524 vss.n102 vss.n101 42250
R1525 vss.n98 vss.n97 42250
R1526 vss.n94 vss.n93 42250
R1527 vss.n90 vss.n89 42250
R1528 vss.n86 vss.n1 40867.3
R1529 vss.n87 vss.n86 13561.1
R1530 vss.n119 vss.n118 13560.9
R1531 vss.n115 vss.n114 13560.9
R1532 vss.n111 vss.n110 13560.9
R1533 vss.n107 vss.n106 13560.9
R1534 vss.n103 vss.n102 13560.9
R1535 vss.n99 vss.n98 13560.9
R1536 vss.n95 vss.n94 13560.9
R1537 vss.n91 vss.n90 13560.9
R1538 vss.n118 vss.n77 4104.97
R1539 vss.n114 vss.n78 4104.97
R1540 vss.n110 vss.n79 4104.97
R1541 vss.n106 vss.n80 4104.97
R1542 vss.n102 vss.n81 4104.97
R1543 vss.n98 vss.n82 4104.97
R1544 vss.n94 vss.n83 4104.97
R1545 vss.n90 vss.n84 4104.97
R1546 vss.n86 vss.n85 3523.68
R1547 vss.t177 vss.t179 1631.65
R1548 vss.t151 vss.t110 1631.65
R1549 vss.t132 vss.t134 1611.86
R1550 vss.t302 vss.t292 1611.86
R1551 vss.t369 vss.t367 1611.86
R1552 vss.t97 vss.t188 1611.86
R1553 vss.t120 vss.t118 1611.86
R1554 vss.t29 vss.t56 1611.86
R1555 vss.t378 vss.t380 1611.86
R1556 vss.t107 vss.t271 1611.86
R1557 vss.t142 vss.t140 1611.86
R1558 vss.t258 vss.t255 1611.86
R1559 vss.t327 vss.t329 1611.86
R1560 vss.t123 vss.t374 1611.86
R1561 vss.t361 vss.t363 1611.86
R1562 vss.t163 vss.t32 1611.86
R1563 vss.t336 vss.t338 1611.86
R1564 vss.t273 vss.t228 1611.86
R1565 vss.t86 vss.t84 1611.86
R1566 vss.t146 vss.t284 1611.86
R1567 vss.n2 vss.t112 1294.68
R1568 vss.t278 vss.n74 1278.98
R1569 vss.t93 vss.n66 1278.98
R1570 vss.t8 vss.n58 1278.98
R1571 vss.t266 vss.n50 1278.98
R1572 vss.t253 vss.n42 1278.98
R1573 vss.t357 vss.n34 1278.98
R1574 vss.t406 vss.n26 1278.98
R1575 vss.t316 vss.n18 1278.98
R1576 vss.t344 vss.n10 1278.98
R1577 vss.t4 vss.t109 1152.8
R1578 vss.t110 vss.t193 1152.8
R1579 vss vss.t181 1148.36
R1580 vss.t125 vss.t291 1138.81
R1581 vss.t292 vss.t191 1138.81
R1582 vss.t221 vss.t190 1138.81
R1583 vss.t188 vss.t219 1138.81
R1584 vss.t376 vss.t55 1138.81
R1585 vss.t56 vss.t400 1138.81
R1586 vss.t153 vss.t270 1138.81
R1587 vss.t271 vss.t195 1138.81
R1588 vss.t350 vss.t257 1138.81
R1589 vss.t255 vss.t36 1138.81
R1590 vss.t90 vss.t373 1138.81
R1591 vss.t374 vss.t404 1138.81
R1592 vss.t116 vss.t31 1138.81
R1593 vss.t32 vss.t34 1138.81
R1594 vss.t275 vss.t230 1138.81
R1595 vss.t228 vss.t217 1138.81
R1596 vss.t148 vss.t286 1138.81
R1597 vss.t284 vss.t402 1138.81
R1598 vss vss.t205 1134.43
R1599 vss vss.t206 1134.43
R1600 vss vss.t41 1134.43
R1601 vss vss.t182 1134.43
R1602 vss vss.t0 1134.43
R1603 vss vss.t1 1134.43
R1604 vss vss.t42 1134.43
R1605 vss vss.t63 1134.43
R1606 vss vss.t184 1134.43
R1607 vss vss.t177 1117.33
R1608 vss vss.t132 1103.77
R1609 vss vss.t369 1103.77
R1610 vss vss.t120 1103.77
R1611 vss vss.t378 1103.77
R1612 vss vss.t142 1103.77
R1613 vss vss.t327 1103.77
R1614 vss vss.t361 1103.77
R1615 vss vss.t336 1103.77
R1616 vss vss.t86 1103.77
R1617 vss.t179 vss.t4 993.179
R1618 vss.t109 vss.t131 993.179
R1619 vss.t134 vss.t125 981.133
R1620 vss.t291 vss.t64 981.133
R1621 vss.t367 vss.t221 981.133
R1622 vss.t190 vss.t249 981.133
R1623 vss.t118 vss.t376 981.133
R1624 vss.t55 vss.t136 981.133
R1625 vss.t380 vss.t153 981.133
R1626 vss.t270 vss.t38 981.133
R1627 vss.t140 vss.t350 981.133
R1628 vss.t257 vss.t150 981.133
R1629 vss.t329 vss.t90 981.133
R1630 vss.t373 vss.t162 981.133
R1631 vss.t363 vss.t116 981.133
R1632 vss.t31 vss.t277 981.133
R1633 vss.t338 vss.t275 981.133
R1634 vss.t230 vss.t122 981.133
R1635 vss.t84 vss.t148 981.133
R1636 vss.t286 vss.t145 981.133
R1637 vss.t181 vss.t80 815.826
R1638 vss vss.n2 815.826
R1639 vss.t205 vss.t334 805.931
R1640 vss vss.n74 805.931
R1641 vss.t206 vss.t325 805.931
R1642 vss vss.n66 805.931
R1643 vss.t41 vss.t167 805.931
R1644 vss vss.n58 805.931
R1645 vss.t182 vss.t352 805.931
R1646 vss vss.n50 805.931
R1647 vss.t0 vss.t173 805.931
R1648 vss vss.n42 805.931
R1649 vss.t1 vss.t127 805.931
R1650 vss vss.n34 805.931
R1651 vss.t42 vss.t314 805.931
R1652 vss vss.n26 805.931
R1653 vss.t63 vss.t158 805.931
R1654 vss vss.n18 805.931
R1655 vss.t184 vss.t346 805.931
R1656 vss vss.n10 805.931
R1657 vss.n70 vss.n69 805.874
R1658 vss.n62 vss.n61 805.874
R1659 vss.n54 vss.n53 805.874
R1660 vss.n46 vss.n45 805.874
R1661 vss.n38 vss.n37 805.874
R1662 vss.n30 vss.n29 805.874
R1663 vss.n22 vss.n21 805.874
R1664 vss.n14 vss.n13 805.874
R1665 vss.n6 vss.n5 805.874
R1666 vss.n77 vss.t243 760.808
R1667 vss.n78 vss.t82 760.808
R1668 vss.n79 vss.t226 760.808
R1669 vss.n80 vss.t58 760.808
R1670 vss.n81 vss.t6 760.808
R1671 vss.n82 vss.t39 760.808
R1672 vss.n83 vss.t88 760.808
R1673 vss.n84 vss.t215 760.808
R1674 vss.t131 vss.t151 744.885
R1675 vss.t64 vss.t302 735.85
R1676 vss.t249 vss.t97 735.85
R1677 vss.t136 vss.t29 735.85
R1678 vss.t38 vss.t107 735.85
R1679 vss.t150 vss.t258 735.85
R1680 vss.t162 vss.t123 735.85
R1681 vss.t277 vss.t163 735.85
R1682 vss.t122 vss.t273 735.85
R1683 vss.t145 vss.t146 735.85
R1684 vss.t112 vss.n1 696.112
R1685 vss.n85 vss.t365 638.866
R1686 vss.t27 vss.t233 593.802
R1687 vss.t308 vss.t237 593.802
R1688 vss.t207 vss.t247 593.802
R1689 vss.t49 vss.t231 593.802
R1690 vss.t69 vss.t239 593.802
R1691 vss.t15 vss.t262 593.802
R1692 vss.t382 vss.t264 593.802
R1693 vss.t104 vss.t235 593.802
R1694 vss.t299 vss.t260 593.802
R1695 vss.t80 vss 518.759
R1696 vss.t193 vss 514.326
R1697 vss.t334 vss 512.466
R1698 vss.t325 vss 512.466
R1699 vss.t167 vss 512.466
R1700 vss.t352 vss 512.466
R1701 vss.t173 vss 512.466
R1702 vss.t127 vss 512.466
R1703 vss.t314 vss 512.466
R1704 vss.t158 vss 512.466
R1705 vss.t346 vss 512.466
R1706 vss.t393 vss 508.087
R1707 vss.t191 vss 508.087
R1708 vss.t243 vss 508.087
R1709 vss.t219 vss 508.087
R1710 vss.t82 vss 508.087
R1711 vss.t400 vss 508.087
R1712 vss.t226 vss 508.087
R1713 vss.t195 vss 508.087
R1714 vss.t58 vss 508.087
R1715 vss.t36 vss 508.087
R1716 vss.t6 vss 508.087
R1717 vss.t404 vss 508.087
R1718 vss.t39 vss 508.087
R1719 vss.t34 vss 508.087
R1720 vss.t88 vss 508.087
R1721 vss.t217 vss 508.087
R1722 vss.t215 vss 508.087
R1723 vss.t402 vss 508.087
R1724 vss vss.n0 467.339
R1725 vss.n119 vss 408.238
R1726 vss.n115 vss 408.238
R1727 vss.n111 vss 408.238
R1728 vss.n107 vss 408.238
R1729 vss.n103 vss 408.238
R1730 vss.n99 vss 408.238
R1731 vss.n95 vss 408.238
R1732 vss.n91 vss 408.238
R1733 vss.n87 vss 408.238
R1734 vss.n283 vss.t60 381.882
R1735 vss.t203 vss.t241 355.178
R1736 vss.t365 vss 352.079
R1737 vss.n120 vss.t280 349.329
R1738 vss.n116 vss.t95 349.329
R1739 vss.n112 vss.t10 349.329
R1740 vss.n108 vss.t268 349.329
R1741 vss.n104 vss.t251 349.329
R1742 vss.n100 vss.t359 349.329
R1743 vss.n96 vss.t408 349.329
R1744 vss.n92 vss.t318 349.329
R1745 vss.n88 vss.t342 349.329
R1746 vss.n85 vss.n5 347.269
R1747 vss vss.t203 309.779
R1748 vss.t241 vss 309.779
R1749 vss.t233 vss 307.505
R1750 vss.t237 vss 307.505
R1751 vss.t247 vss 307.505
R1752 vss.t231 vss 307.505
R1753 vss.t239 vss 307.505
R1754 vss.t262 vss 307.505
R1755 vss.t264 vss 307.505
R1756 vss.t235 vss 307.505
R1757 vss.t260 vss 307.505
R1758 vss.n121 vss.t278 289.084
R1759 vss.n117 vss.t93 289.084
R1760 vss.n113 vss.t8 289.084
R1761 vss.n109 vss.t266 289.084
R1762 vss.n105 vss.t253 289.084
R1763 vss.n101 vss.t357 289.084
R1764 vss.n97 vss.t406 289.084
R1765 vss.n93 vss.t316 289.084
R1766 vss.n89 vss.t344 289.084
R1767 vss.n283 vss.t199 286.949
R1768 vss.n71 vss.n70 265.091
R1769 vss.n63 vss.n62 265.091
R1770 vss.n55 vss.n54 265.091
R1771 vss.n47 vss.n46 265.091
R1772 vss.n39 vss.n38 265.091
R1773 vss.n31 vss.n30 265.091
R1774 vss.n23 vss.n22 265.091
R1775 vss.n15 vss.n14 265.091
R1776 vss.n7 vss.n6 265.091
R1777 vss.t21 vss.t23 249.52
R1778 vss.t22 vss.t24 249.52
R1779 vss.t310 vss.t306 249.52
R1780 vss.t311 vss.t304 249.52
R1781 vss.t210 vss.t211 249.52
R1782 vss.t214 vss.t209 249.52
R1783 vss.t53 vss.t54 249.52
R1784 vss.t51 vss.t52 249.52
R1785 vss.t71 vss.t73 249.52
R1786 vss.t72 vss.t74 249.52
R1787 vss.t18 vss.t12 249.52
R1788 vss.t19 vss.t17 249.52
R1789 vss.t388 vss.t384 249.52
R1790 vss.t389 vss.t385 249.52
R1791 vss.t101 vss.t99 249.52
R1792 vss.t106 vss.t100 249.52
R1793 vss.t301 vss.t296 249.52
R1794 vss.t294 vss.t295 249.52
R1795 vss.t200 vss.t197 249.52
R1796 vss.n77 vss.n69 225.327
R1797 vss.n78 vss.n61 225.327
R1798 vss.n79 vss.n53 225.327
R1799 vss.n80 vss.n45 225.327
R1800 vss.n81 vss.n37 225.327
R1801 vss.n82 vss.n29 225.327
R1802 vss.n83 vss.n21 225.327
R1803 vss.n84 vss.n13 225.327
R1804 vss vss.n71 222.675
R1805 vss vss.n63 222.675
R1806 vss vss.n55 222.675
R1807 vss vss.n47 222.675
R1808 vss vss.n39 222.675
R1809 vss vss.n31 222.675
R1810 vss vss.n23 222.675
R1811 vss vss.n15 222.675
R1812 vss vss.n7 222.675
R1813 vss.t26 vss.t390 215.212
R1814 vss.t307 vss.t287 215.212
R1815 vss.t212 vss.t185 215.212
R1816 vss.t47 vss.t223 215.212
R1817 vss.t68 vss.t137 215.212
R1818 vss.t14 vss.t397 215.212
R1819 vss.t386 vss.t157 215.212
R1820 vss.t102 vss.t75 215.212
R1821 vss.t297 vss.t43 215.212
R1822 vss vss.t391 212.072
R1823 vss vss.t288 212.072
R1824 vss vss.t186 212.072
R1825 vss vss.t224 212.072
R1826 vss vss.t138 212.072
R1827 vss vss.t395 212.072
R1828 vss vss.t155 212.072
R1829 vss vss.t76 212.072
R1830 vss vss.t44 212.072
R1831 vss.t323 vss.n119 208.974
R1832 vss.t165 vss.n115 208.974
R1833 vss.t354 vss.n111 208.974
R1834 vss.t171 vss.n107 208.974
R1835 vss.t129 vss.n103 208.974
R1836 vss.t312 vss.n99 208.974
R1837 vss.t160 vss.n95 208.974
R1838 vss.t348 vss.n91 208.974
R1839 vss.t78 vss.n87 208.974
R1840 vss.t114 vss.n282 207.415
R1841 vss.t340 vss.t26 190.26
R1842 vss.t398 vss.t307 190.26
R1843 vss.t282 vss.t212 190.26
R1844 vss.t320 vss.t47 190.26
R1845 vss.t169 vss.t68 190.26
R1846 vss.t371 vss.t14 190.26
R1847 vss.t175 vss.t386 190.26
R1848 vss.t65 vss.t102 190.26
R1849 vss.t332 vss.t297 190.26
R1850 vss.t245 vss.t198 185.582
R1851 vss.t322 vss.t25 184.022
R1852 vss.t331 vss.t305 184.022
R1853 vss.t46 vss.t213 184.022
R1854 vss.t250 vss.t48 184.022
R1855 vss.t92 vss.t67 184.022
R1856 vss.t144 vss.t13 184.022
R1857 vss.t290 vss.t387 184.022
R1858 vss.t183 vss.t103 184.022
R1859 vss.t356 vss.t298 184.022
R1860 vss.t201 vss.t114 182.463
R1861 vss.t202 vss.t62 176.225
R1862 vss.t20 vss.t202 173.106
R1863 vss.t2 vss.t201 166.868
R1864 vss.n121 vss.n120 121.641
R1865 vss.n117 vss.n116 121.641
R1866 vss.n113 vss.n112 121.641
R1867 vss.n109 vss.n108 121.641
R1868 vss.n105 vss.n104 121.641
R1869 vss.n101 vss.n100 121.641
R1870 vss.n97 vss.n96 121.641
R1871 vss.n93 vss.n92 121.641
R1872 vss.n89 vss.n88 121.641
R1873 vss.n282 vss.n1 121.641
R1874 vss.t391 vss.t27 95.4328
R1875 vss.t288 vss.t308 95.4328
R1876 vss.t186 vss.t207 95.4328
R1877 vss.t224 vss.t49 95.4328
R1878 vss.t138 vss.t69 95.4328
R1879 vss.t395 vss.t15 95.4328
R1880 vss.t155 vss.t382 95.4328
R1881 vss.t76 vss.t104 95.4328
R1882 vss.t44 vss.t299 95.4328
R1883 vss.t197 vss.t2 82.6541
R1884 vss.t25 vss.t323 77.9755
R1885 vss.t305 vss.t165 77.9755
R1886 vss.t213 vss.t354 77.9755
R1887 vss.t48 vss.t171 77.9755
R1888 vss.t67 vss.t129 77.9755
R1889 vss.t13 vss.t312 77.9755
R1890 vss.t387 vss.t160 77.9755
R1891 vss.t103 vss.t348 77.9755
R1892 vss.t298 vss.t78 77.9755
R1893 vss.t198 vss.t20 76.4161
R1894 vss.t62 vss.t200 73.297
R1895 vss.n122 vss.t393 72.5527
R1896 vss.t24 vss.t322 65.4995
R1897 vss.t304 vss.t331 65.4995
R1898 vss.t209 vss.t46 65.4995
R1899 vss.t52 vss.t250 65.4995
R1900 vss.t74 vss.t92 65.4995
R1901 vss.t17 vss.t144 65.4995
R1902 vss.t385 vss.t290 65.4995
R1903 vss.t100 vss.t183 65.4995
R1904 vss.t295 vss.t356 65.4995
R1905 vss.t199 vss.t245 63.94
R1906 vss.t23 vss.t340 59.2615
R1907 vss.t306 vss.t398 59.2615
R1908 vss.t211 vss.t282 59.2615
R1909 vss.t54 vss.t320 59.2615
R1910 vss.t73 vss.t169 59.2615
R1911 vss.t12 vss.t371 59.2615
R1912 vss.t384 vss.t175 59.2615
R1913 vss.t99 vss.t65 59.2615
R1914 vss.t296 vss.t332 59.2615
R1915 vss.t280 vss.t21 40.5475
R1916 vss.t95 vss.t310 40.5475
R1917 vss.t10 vss.t210 40.5475
R1918 vss.t268 vss.t53 40.5475
R1919 vss.t251 vss.t71 40.5475
R1920 vss.t359 vss.t18 40.5475
R1921 vss.t408 vss.t388 40.5475
R1922 vss.t318 vss.t101 40.5475
R1923 vss.t342 vss.t301 40.5475
R1924 vss.t390 vss.t22 34.3095
R1925 vss.t287 vss.t311 34.3095
R1926 vss.t185 vss.t214 34.3095
R1927 vss.t223 vss.t51 34.3095
R1928 vss.t137 vss.t72 34.3095
R1929 vss.t397 vss.t19 34.3095
R1930 vss.t157 vss.t389 34.3095
R1931 vss.t75 vss.t106 34.3095
R1932 vss.t43 vss.t294 34.3095
R1933 vss.t60 vss 29.376
R1934 vss.n284 vss.n0 24.035
R1935 vss.n279 vss.t246 8.79702
R1936 vss.n271 vss.t152 8.79702
R1937 vss.n261 vss.t79 8.79702
R1938 vss.n255 vss.t147 8.79702
R1939 vss.n245 vss.t349 8.79702
R1940 vss.n239 vss.t274 8.79702
R1941 vss.n229 vss.t161 8.79702
R1942 vss.n223 vss.t164 8.79702
R1943 vss.n213 vss.t313 8.79702
R1944 vss.n207 vss.t124 8.79702
R1945 vss.n197 vss.t130 8.79702
R1946 vss.n191 vss.t259 8.79702
R1947 vss.n181 vss.t172 8.79702
R1948 vss.n175 vss.t108 8.79702
R1949 vss.n165 vss.t355 8.79702
R1950 vss.n159 vss.t30 8.79702
R1951 vss.n149 vss.t166 8.79702
R1952 vss.n143 vss.t98 8.79702
R1953 vss.n133 vss.t324 8.79702
R1954 vss.n127 vss.t303 8.79702
R1955 vss.n277 vss.n276 6.40811
R1956 vss.n272 vss.n3 6.40811
R1957 vss.n263 vss.n8 6.40811
R1958 vss.n256 vss.n11 6.40811
R1959 vss.n247 vss.n16 6.40811
R1960 vss.n240 vss.n19 6.40811
R1961 vss.n231 vss.n24 6.40811
R1962 vss.n224 vss.n27 6.40811
R1963 vss.n215 vss.n32 6.40811
R1964 vss.n208 vss.n35 6.40811
R1965 vss.n199 vss.n40 6.40811
R1966 vss.n192 vss.n43 6.40811
R1967 vss.n183 vss.n48 6.40811
R1968 vss.n176 vss.n51 6.40811
R1969 vss.n167 vss.n56 6.40811
R1970 vss.n160 vss.n59 6.40811
R1971 vss.n151 vss.n64 6.40811
R1972 vss.n144 vss.n67 6.40811
R1973 vss.n135 vss.n72 6.40811
R1974 vss.n128 vss.n75 6.40811
R1975 vss.n270 vss.n4 6.4042
R1976 vss.n280 vss.n275 6.4042
R1977 vss.n254 vss.n12 6.4042
R1978 vss.n260 vss.n9 6.4042
R1979 vss.n238 vss.n20 6.4042
R1980 vss.n244 vss.n17 6.4042
R1981 vss.n222 vss.n28 6.4042
R1982 vss.n228 vss.n25 6.4042
R1983 vss.n206 vss.n36 6.4042
R1984 vss.n212 vss.n33 6.4042
R1985 vss.n190 vss.n44 6.4042
R1986 vss.n196 vss.n41 6.4042
R1987 vss.n174 vss.n52 6.4042
R1988 vss.n180 vss.n49 6.4042
R1989 vss.n158 vss.n60 6.4042
R1990 vss.n164 vss.n57 6.4042
R1991 vss.n142 vss.n68 6.4042
R1992 vss.n148 vss.n65 6.4042
R1993 vss.n126 vss.n76 6.4042
R1994 vss.n132 vss.n73 6.4042
R1995 vss.n264 vss.n7 5.28469
R1996 vss.n248 vss.n15 5.28469
R1997 vss.n232 vss.n23 5.28469
R1998 vss.n216 vss.n31 5.28469
R1999 vss.n200 vss.n39 5.28469
R2000 vss.n184 vss.n47 5.28469
R2001 vss.n168 vss.n55 5.28469
R2002 vss.n152 vss.n63 5.28469
R2003 vss.n136 vss.n71 5.28469
R2004 vss.n286 vss.n0 5.28469
R2005 vss.n267 vss.t366 4.63989
R2006 vss.n269 vss.t178 4.63989
R2007 vss.n274 vss.t113 4.63989
R2008 vss.n262 vss.t300 4.63989
R2009 vss.n251 vss.t216 4.63989
R2010 vss.n253 vss.t87 4.63989
R2011 vss.n258 vss.t345 4.63989
R2012 vss.n246 vss.t105 4.63989
R2013 vss.n235 vss.t89 4.63989
R2014 vss.n237 vss.t337 4.63989
R2015 vss.n242 vss.t317 4.63989
R2016 vss.n230 vss.t383 4.63989
R2017 vss.n219 vss.t40 4.63989
R2018 vss.n221 vss.t362 4.63989
R2019 vss.n226 vss.t407 4.63989
R2020 vss.n214 vss.t16 4.63989
R2021 vss.n203 vss.t7 4.63989
R2022 vss.n205 vss.t328 4.63989
R2023 vss.n210 vss.t358 4.63989
R2024 vss.n198 vss.t70 4.63989
R2025 vss.n187 vss.t59 4.63989
R2026 vss.n189 vss.t143 4.63989
R2027 vss.n194 vss.t254 4.63989
R2028 vss.n182 vss.t50 4.63989
R2029 vss.n171 vss.t227 4.63989
R2030 vss.n173 vss.t379 4.63989
R2031 vss.n178 vss.t267 4.63989
R2032 vss.n166 vss.t208 4.63989
R2033 vss.n155 vss.t83 4.63989
R2034 vss.n157 vss.t121 4.63989
R2035 vss.n162 vss.t9 4.63989
R2036 vss.n150 vss.t309 4.63989
R2037 vss.n139 vss.t244 4.63989
R2038 vss.n141 vss.t370 4.63989
R2039 vss.n146 vss.t94 4.63989
R2040 vss.n134 vss.t28 4.63989
R2041 vss.n123 vss.t394 4.63989
R2042 vss.n125 vss.t133 4.63989
R2043 vss.n130 vss.t279 4.63989
R2044 vss.n278 vss.t204 4.63989
R2045 vss.n268 vss.t81 4.51271
R2046 vss.n252 vss.t347 4.51271
R2047 vss.n236 vss.t159 4.51271
R2048 vss.n220 vss.t315 4.51271
R2049 vss.n204 vss.t128 4.51271
R2050 vss.n188 vss.t174 4.51271
R2051 vss.n172 vss.t353 4.51271
R2052 vss.n156 vss.t168 4.51271
R2053 vss.n140 vss.t326 4.51271
R2054 vss.n124 vss.t335 4.51271
R2055 vss.n276 vss.t61 3.9605
R2056 vss.n3 vss.t111 3.9605
R2057 vss.n8 vss.t45 3.9605
R2058 vss.n11 vss.t285 3.9605
R2059 vss.n16 vss.t77 3.9605
R2060 vss.n19 vss.t229 3.9605
R2061 vss.n24 vss.t156 3.9605
R2062 vss.n27 vss.t33 3.9605
R2063 vss.n32 vss.t396 3.9605
R2064 vss.n35 vss.t375 3.9605
R2065 vss.n40 vss.t139 3.9605
R2066 vss.n43 vss.t256 3.9605
R2067 vss.n48 vss.t225 3.9605
R2068 vss.n51 vss.t272 3.9605
R2069 vss.n56 vss.t187 3.9605
R2070 vss.n59 vss.t57 3.9605
R2071 vss.n64 vss.t289 3.9605
R2072 vss.n67 vss.t189 3.9605
R2073 vss.n72 vss.t392 3.9605
R2074 vss.n75 vss.t293 3.9605
R2075 vss.n285 vss.n284 3.6294
R2076 vss.n266 vss.n5 3.6294
R2077 vss.n273 vss.n2 3.6294
R2078 vss.n265 vss.n6 3.6294
R2079 vss.n250 vss.n13 3.6294
R2080 vss.n257 vss.n10 3.6294
R2081 vss.n249 vss.n14 3.6294
R2082 vss.n234 vss.n21 3.6294
R2083 vss.n241 vss.n18 3.6294
R2084 vss.n233 vss.n22 3.6294
R2085 vss.n218 vss.n29 3.6294
R2086 vss.n225 vss.n26 3.6294
R2087 vss.n217 vss.n30 3.6294
R2088 vss.n202 vss.n37 3.6294
R2089 vss.n209 vss.n34 3.6294
R2090 vss.n201 vss.n38 3.6294
R2091 vss.n186 vss.n45 3.6294
R2092 vss.n193 vss.n42 3.6294
R2093 vss.n185 vss.n46 3.6294
R2094 vss.n170 vss.n53 3.6294
R2095 vss.n177 vss.n50 3.6294
R2096 vss.n169 vss.n54 3.6294
R2097 vss.n154 vss.n61 3.6294
R2098 vss.n161 vss.n58 3.6294
R2099 vss.n153 vss.n62 3.6294
R2100 vss.n138 vss.n69 3.6294
R2101 vss.n145 vss.n66 3.6294
R2102 vss.n137 vss.n70 3.6294
R2103 vss.n129 vss.n74 3.6294
R2104 vss.n4 vss.t180 2.07392
R2105 vss.n4 vss.t5 2.07392
R2106 vss.n275 vss.t115 2.07392
R2107 vss.n275 vss.t3 2.07392
R2108 vss.n12 vss.t85 2.07392
R2109 vss.n12 vss.t149 2.07392
R2110 vss.n9 vss.t343 2.07392
R2111 vss.n9 vss.t333 2.07392
R2112 vss.n20 vss.t339 2.07392
R2113 vss.n20 vss.t276 2.07392
R2114 vss.n17 vss.t319 2.07392
R2115 vss.n17 vss.t66 2.07392
R2116 vss.n28 vss.t364 2.07392
R2117 vss.n28 vss.t117 2.07392
R2118 vss.n25 vss.t409 2.07392
R2119 vss.n25 vss.t176 2.07392
R2120 vss.n36 vss.t330 2.07392
R2121 vss.n36 vss.t91 2.07392
R2122 vss.n33 vss.t360 2.07392
R2123 vss.n33 vss.t372 2.07392
R2124 vss.n44 vss.t141 2.07392
R2125 vss.n44 vss.t351 2.07392
R2126 vss.n41 vss.t252 2.07392
R2127 vss.n41 vss.t170 2.07392
R2128 vss.n52 vss.t381 2.07392
R2129 vss.n52 vss.t154 2.07392
R2130 vss.n49 vss.t269 2.07392
R2131 vss.n49 vss.t321 2.07392
R2132 vss.n60 vss.t119 2.07392
R2133 vss.n60 vss.t377 2.07392
R2134 vss.n57 vss.t11 2.07392
R2135 vss.n57 vss.t283 2.07392
R2136 vss.n68 vss.t368 2.07392
R2137 vss.n68 vss.t222 2.07392
R2138 vss.n65 vss.t96 2.07392
R2139 vss.n65 vss.t399 2.07392
R2140 vss.n76 vss.t135 2.07392
R2141 vss.n76 vss.t126 2.07392
R2142 vss.n73 vss.t281 2.07392
R2143 vss.n73 vss.t341 2.07392
R2144 vss.n276 vss.t242 1.84987
R2145 vss.n3 vss.t194 1.84987
R2146 vss.n8 vss.t261 1.84987
R2147 vss.n11 vss.t403 1.84987
R2148 vss.n16 vss.t236 1.84987
R2149 vss.n19 vss.t218 1.84987
R2150 vss.n24 vss.t265 1.84987
R2151 vss.n27 vss.t35 1.84987
R2152 vss.n32 vss.t263 1.84987
R2153 vss.n35 vss.t405 1.84987
R2154 vss.n40 vss.t240 1.84987
R2155 vss.n43 vss.t37 1.84987
R2156 vss.n48 vss.t232 1.84987
R2157 vss.n51 vss.t196 1.84987
R2158 vss.n56 vss.t248 1.84987
R2159 vss.n59 vss.t401 1.84987
R2160 vss.n64 vss.t238 1.84987
R2161 vss.n67 vss.t220 1.84987
R2162 vss.n72 vss.t234 1.84987
R2163 vss.n75 vss.t192 1.84987
R2164 vss.n120 vss 1.48621
R2165 vss.n116 vss 1.48621
R2166 vss.n112 vss 1.48621
R2167 vss.n108 vss 1.48621
R2168 vss.n104 vss 1.48621
R2169 vss.n100 vss 1.48621
R2170 vss.n96 vss 1.48621
R2171 vss.n92 vss 1.48621
R2172 vss.n88 vss 1.48621
R2173 vss.n282 vss 1.48621
R2174 vss.n259 vss 0.7205
R2175 vss.n243 vss 0.7205
R2176 vss.n227 vss 0.7205
R2177 vss.n211 vss 0.7205
R2178 vss.n195 vss 0.7205
R2179 vss.n179 vss 0.7205
R2180 vss.n163 vss 0.7205
R2181 vss.n147 vss 0.7205
R2182 vss.n131 vss 0.7205
R2183 vss vss.n281 0.709842
R2184 vss.n270 vss.n269 0.172371
R2185 vss.n254 vss.n253 0.172371
R2186 vss.n238 vss.n237 0.172371
R2187 vss.n222 vss.n221 0.172371
R2188 vss.n206 vss.n205 0.172371
R2189 vss.n190 vss.n189 0.172371
R2190 vss.n174 vss.n173 0.172371
R2191 vss.n158 vss.n157 0.172371
R2192 vss.n142 vss.n141 0.172371
R2193 vss.n126 vss.n125 0.172371
R2194 vss vss.n270 0.132887
R2195 vss.n280 vss 0.132887
R2196 vss vss.n254 0.132887
R2197 vss vss.n260 0.132887
R2198 vss vss.n238 0.132887
R2199 vss vss.n244 0.132887
R2200 vss vss.n222 0.132887
R2201 vss vss.n228 0.132887
R2202 vss vss.n206 0.132887
R2203 vss vss.n212 0.132887
R2204 vss vss.n190 0.132887
R2205 vss vss.n196 0.132887
R2206 vss vss.n174 0.132887
R2207 vss vss.n180 0.132887
R2208 vss vss.n158 0.132887
R2209 vss vss.n164 0.132887
R2210 vss vss.n142 0.132887
R2211 vss vss.n148 0.132887
R2212 vss vss.n126 0.132887
R2213 vss vss.n132 0.132887
R2214 vss.n271 vss 0.122435
R2215 vss.n255 vss 0.122435
R2216 vss.n239 vss 0.122435
R2217 vss.n223 vss 0.122435
R2218 vss.n207 vss 0.122435
R2219 vss.n191 vss 0.122435
R2220 vss.n175 vss 0.122435
R2221 vss.n159 vss 0.122435
R2222 vss.n143 vss 0.122435
R2223 vss.n127 vss 0.122435
R2224 vss vss.n279 0.122412
R2225 vss.n261 vss 0.121383
R2226 vss.n245 vss 0.121383
R2227 vss.n229 vss 0.121383
R2228 vss.n213 vss 0.121383
R2229 vss.n197 vss 0.121383
R2230 vss.n181 vss 0.121383
R2231 vss.n165 vss 0.121383
R2232 vss.n149 vss 0.121383
R2233 vss.n133 vss 0.121383
R2234 vss vss.n272 0.118952
R2235 vss vss.n256 0.118952
R2236 vss vss.n240 0.118952
R2237 vss vss.n224 0.118952
R2238 vss vss.n208 0.118952
R2239 vss vss.n192 0.118952
R2240 vss vss.n176 0.118952
R2241 vss vss.n160 0.118952
R2242 vss vss.n144 0.118952
R2243 vss vss.n128 0.118952
R2244 vss.n272 vss.n271 0.11779
R2245 vss.n256 vss.n255 0.11779
R2246 vss.n240 vss.n239 0.11779
R2247 vss.n224 vss.n223 0.11779
R2248 vss.n208 vss.n207 0.11779
R2249 vss.n192 vss.n191 0.11779
R2250 vss.n176 vss.n175 0.11779
R2251 vss.n160 vss.n159 0.11779
R2252 vss.n144 vss.n143 0.11779
R2253 vss.n128 vss.n127 0.11779
R2254 vss vss.n267 0.102694
R2255 vss vss.n251 0.102694
R2256 vss vss.n235 0.102694
R2257 vss vss.n219 0.102694
R2258 vss vss.n203 0.102694
R2259 vss vss.n187 0.102694
R2260 vss vss.n171 0.102694
R2261 vss vss.n155 0.102694
R2262 vss vss.n139 0.102694
R2263 vss vss.n123 0.102694
R2264 vss.n281 vss.n274 0.101242
R2265 vss.n260 vss.n259 0.0980484
R2266 vss.n244 vss.n243 0.0980484
R2267 vss.n228 vss.n227 0.0980484
R2268 vss.n212 vss.n211 0.0980484
R2269 vss.n196 vss.n195 0.0980484
R2270 vss.n180 vss.n179 0.0980484
R2271 vss.n164 vss.n163 0.0980484
R2272 vss.n148 vss.n147 0.0980484
R2273 vss.n132 vss.n131 0.0980484
R2274 vss vss.n266 0.0957258
R2275 vss vss.n250 0.0957258
R2276 vss vss.n234 0.0957258
R2277 vss vss.n218 0.0957258
R2278 vss vss.n202 0.0957258
R2279 vss vss.n186 0.0957258
R2280 vss vss.n170 0.0957258
R2281 vss vss.n154 0.0957258
R2282 vss vss.n138 0.0957258
R2283 vss vss.n122 0.0957258
R2284 vss.n259 vss.n258 0.0748226
R2285 vss.n243 vss.n242 0.0748226
R2286 vss.n227 vss.n226 0.0748226
R2287 vss.n211 vss.n210 0.0748226
R2288 vss.n195 vss.n194 0.0748226
R2289 vss.n179 vss.n178 0.0748226
R2290 vss.n163 vss.n162 0.0748226
R2291 vss.n147 vss.n146 0.0748226
R2292 vss.n131 vss.n130 0.0748226
R2293 vss.n281 vss.n280 0.071629
R2294 vss.n279 vss.n278 0.071286
R2295 vss.n268 vss 0.0605968
R2296 vss.n252 vss 0.0605968
R2297 vss.n236 vss 0.0605968
R2298 vss.n220 vss 0.0605968
R2299 vss.n204 vss 0.0605968
R2300 vss.n188 vss 0.0605968
R2301 vss.n172 vss 0.0605968
R2302 vss.n156 vss 0.0605968
R2303 vss.n140 vss 0.0605968
R2304 vss.n124 vss 0.0605968
R2305 vss.n274 vss.n273 0.0515968
R2306 vss.n258 vss.n257 0.0515968
R2307 vss.n242 vss.n241 0.0515968
R2308 vss.n226 vss.n225 0.0515968
R2309 vss.n210 vss.n209 0.0515968
R2310 vss.n194 vss.n193 0.0515968
R2311 vss.n178 vss.n177 0.0515968
R2312 vss.n162 vss.n161 0.0515968
R2313 vss.n146 vss.n145 0.0515968
R2314 vss.n130 vss.n129 0.0515968
R2315 vss.n267 vss 0.044629
R2316 vss.n251 vss 0.044629
R2317 vss.n235 vss 0.044629
R2318 vss.n219 vss 0.044629
R2319 vss.n203 vss 0.044629
R2320 vss.n187 vss 0.044629
R2321 vss.n171 vss 0.044629
R2322 vss.n155 vss 0.044629
R2323 vss.n139 vss 0.044629
R2324 vss.n123 vss 0.044629
R2325 vss.n262 vss.n261 0.043835
R2326 vss.n246 vss.n245 0.043835
R2327 vss.n230 vss.n229 0.043835
R2328 vss.n214 vss.n213 0.043835
R2329 vss.n198 vss.n197 0.043835
R2330 vss.n182 vss.n181 0.043835
R2331 vss.n166 vss.n165 0.043835
R2332 vss.n150 vss.n149 0.043835
R2333 vss.n134 vss.n133 0.043835
R2334 vss.n269 vss.n268 0.0425968
R2335 vss.n253 vss.n252 0.0425968
R2336 vss.n237 vss.n236 0.0425968
R2337 vss.n221 vss.n220 0.0425968
R2338 vss.n205 vss.n204 0.0425968
R2339 vss.n189 vss.n188 0.0425968
R2340 vss.n173 vss.n172 0.0425968
R2341 vss.n157 vss.n156 0.0425968
R2342 vss.n141 vss.n140 0.0425968
R2343 vss.n125 vss.n124 0.0425968
R2344 vss vss.n286 0.0413758
R2345 vss.n264 vss 0.04064
R2346 vss.n248 vss 0.04064
R2347 vss.n232 vss 0.04064
R2348 vss.n216 vss 0.04064
R2349 vss.n200 vss 0.04064
R2350 vss.n184 vss 0.04064
R2351 vss.n168 vss 0.04064
R2352 vss.n152 vss 0.04064
R2353 vss.n136 vss 0.04064
R2354 vss vss.n265 0.0338174
R2355 vss vss.n249 0.0338174
R2356 vss vss.n233 0.0338174
R2357 vss vss.n217 0.0338174
R2358 vss vss.n201 0.0338174
R2359 vss vss.n185 0.0338174
R2360 vss vss.n169 0.0338174
R2361 vss vss.n153 0.0338174
R2362 vss vss.n137 0.0338174
R2363 vss.n285 vss 0.0283615
R2364 vss vss.n262 0.02786
R2365 vss vss.n246 0.02786
R2366 vss vss.n230 0.02786
R2367 vss vss.n214 0.02786
R2368 vss vss.n198 0.02786
R2369 vss vss.n182 0.02786
R2370 vss vss.n166 0.02786
R2371 vss vss.n150 0.02786
R2372 vss vss.n134 0.02786
R2373 vss.n278 vss.n277 0.0248788
R2374 vss vss.n263 0.01634
R2375 vss vss.n247 0.01634
R2376 vss vss.n231 0.01634
R2377 vss vss.n215 0.01634
R2378 vss vss.n199 0.01634
R2379 vss vss.n183 0.01634
R2380 vss vss.n167 0.01634
R2381 vss vss.n151 0.01634
R2382 vss vss.n135 0.01634
R2383 vss.n263 vss 0.01346
R2384 vss.n247 vss 0.01346
R2385 vss.n231 vss 0.01346
R2386 vss.n215 vss 0.01346
R2387 vss.n199 vss 0.01346
R2388 vss.n183 vss 0.01346
R2389 vss.n167 vss 0.01346
R2390 vss.n151 vss 0.01346
R2391 vss.n135 vss 0.01346
R2392 vss.n277 vss 0.00398269
R2393 vss.n266 vss 0.00282258
R2394 vss.n273 vss 0.00282258
R2395 vss.n250 vss 0.00282258
R2396 vss.n257 vss 0.00282258
R2397 vss.n234 vss 0.00282258
R2398 vss.n241 vss 0.00282258
R2399 vss.n218 vss 0.00282258
R2400 vss.n225 vss 0.00282258
R2401 vss.n202 vss 0.00282258
R2402 vss.n209 vss 0.00282258
R2403 vss.n186 vss 0.00282258
R2404 vss.n193 vss 0.00282258
R2405 vss.n170 vss 0.00282258
R2406 vss.n177 vss 0.00282258
R2407 vss.n154 vss 0.00282258
R2408 vss.n161 vss 0.00282258
R2409 vss.n138 vss 0.00282258
R2410 vss.n145 vss 0.00282258
R2411 vss.n122 vss 0.00282258
R2412 vss.n129 vss 0.00282258
R2413 vss vss.n285 0.0019664
R2414 vss.n265 vss 0.00194
R2415 vss.n249 vss 0.00194
R2416 vss.n233 vss 0.00194
R2417 vss.n217 vss 0.00194
R2418 vss.n201 vss 0.00194
R2419 vss.n185 vss 0.00194
R2420 vss.n169 vss 0.00194
R2421 vss.n153 vss 0.00194
R2422 vss.n137 vss 0.00194
R2423 vss.n286 vss 0.0012332
R2424 vss vss.n264 0.00122
R2425 vss vss.n248 0.00122
R2426 vss vss.n232 0.00122
R2427 vss vss.n216 0.00122
R2428 vss vss.n200 0.00122
R2429 vss vss.n184 0.00122
R2430 vss vss.n168 0.00122
R2431 vss vss.n152 0.00122
R2432 vss vss.n136 0.00122
R2433 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.7994
R2434 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R2435 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R2436 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R2437 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R2438 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R2439 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R2440 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R2441 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R2442 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R2443 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R2444 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R2445 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R2446 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2447 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R2448 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R2449 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R2450 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R2451 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R2452 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R2453 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R2454 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R2455 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R2456 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R2457 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R2458 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R2459 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R2460 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R2461 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R2462 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R2463 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R2464 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R2465 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R2466 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R2467 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R2468 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R2469 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R2470 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R2471 BUS[1].n2 BUS[1].n0 15.3751
R2472 BUS[1].n9 BUS[1].n7 15.2168
R2473 BUS[1].n2 BUS[1].n1 15.0151
R2474 BUS[1].n4 BUS[1].n3 15.0151
R2475 BUS[1].n21 BUS[1].n20 14.8568
R2476 BUS[1].n19 BUS[1].n18 14.8568
R2477 BUS[1].n17 BUS[1].n16 14.8568
R2478 BUS[1].n15 BUS[1].n14 14.8568
R2479 BUS[1].n13 BUS[1].n12 14.8568
R2480 BUS[1].n11 BUS[1].n10 14.8568
R2481 BUS[1].n9 BUS[1].n8 14.8568
R2482 BUS[1].n6 BUS[1].n5 14.8568
R2483 BUS[1].n22 BUS[1] 0.927417
R2484 BUS[1].n6 BUS[1].n4 0.8825
R2485 BUS[1].n20 BUS[1].t2 0.4555
R2486 BUS[1].n20 BUS[1].t10 0.4555
R2487 BUS[1].n18 BUS[1].t9 0.4555
R2488 BUS[1].n18 BUS[1].t17 0.4555
R2489 BUS[1].n16 BUS[1].t5 0.4555
R2490 BUS[1].n16 BUS[1].t12 0.4555
R2491 BUS[1].n14 BUS[1].t11 0.4555
R2492 BUS[1].n14 BUS[1].t14 0.4555
R2493 BUS[1].n12 BUS[1].t1 0.4555
R2494 BUS[1].n12 BUS[1].t4 0.4555
R2495 BUS[1].n10 BUS[1].t8 0.4555
R2496 BUS[1].n10 BUS[1].t16 0.4555
R2497 BUS[1].n8 BUS[1].t15 0.4555
R2498 BUS[1].n8 BUS[1].t7 0.4555
R2499 BUS[1].n7 BUS[1].t6 0.4555
R2500 BUS[1].n7 BUS[1].t13 0.4555
R2501 BUS[1].n5 BUS[1].t0 0.4555
R2502 BUS[1].n5 BUS[1].t3 0.4555
R2503 BUS[1].n0 BUS[1].t19 0.41
R2504 BUS[1].n0 BUS[1].t20 0.41
R2505 BUS[1].n1 BUS[1].t21 0.41
R2506 BUS[1].n1 BUS[1].t23 0.41
R2507 BUS[1].n3 BUS[1].t22 0.41
R2508 BUS[1].n3 BUS[1].t18 0.41
R2509 BUS[1].n4 BUS[1].n2 0.3605
R2510 BUS[1].n11 BUS[1].n9 0.3605
R2511 BUS[1].n13 BUS[1].n11 0.3605
R2512 BUS[1].n15 BUS[1].n13 0.3605
R2513 BUS[1].n17 BUS[1].n15 0.3605
R2514 BUS[1].n19 BUS[1].n17 0.3605
R2515 BUS[1].n21 BUS[1].n19 0.3605
R2516 BUS[1].n22 BUS[1].n6 0.203
R2517 BUS[1] BUS[1].n22 0.0430197
R2518 BUS[1].n22 BUS[1].n21 0.015125
R2519 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.7994
R2520 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R2521 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R2522 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R2523 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R2524 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R2525 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R2526 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R2527 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R2528 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R2529 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R2530 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R2531 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R2532 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2533 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R2534 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R2535 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R2536 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R2537 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R2538 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R2539 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R2540 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R2541 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R2542 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R2543 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R2544 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R2545 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R2546 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R2547 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R2548 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R2549 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R2550 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R2551 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R2552 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R2553 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R2554 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R2555 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R2556 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R2557 BUS[5].n2 BUS[5].n0 15.3751
R2558 BUS[5].n9 BUS[5].n7 15.2168
R2559 BUS[5].n2 BUS[5].n1 15.0151
R2560 BUS[5].n4 BUS[5].n3 15.0151
R2561 BUS[5].n21 BUS[5].n20 14.8568
R2562 BUS[5].n19 BUS[5].n18 14.8568
R2563 BUS[5].n17 BUS[5].n16 14.8568
R2564 BUS[5].n15 BUS[5].n14 14.8568
R2565 BUS[5].n13 BUS[5].n12 14.8568
R2566 BUS[5].n11 BUS[5].n10 14.8568
R2567 BUS[5].n9 BUS[5].n8 14.8568
R2568 BUS[5].n6 BUS[5].n5 14.8568
R2569 BUS[5].n22 BUS[5] 0.921051
R2570 BUS[5].n6 BUS[5].n4 0.8825
R2571 BUS[5].n20 BUS[5].t13 0.4555
R2572 BUS[5].n20 BUS[5].t16 0.4555
R2573 BUS[5].n18 BUS[5].t21 0.4555
R2574 BUS[5].n18 BUS[5].t23 0.4555
R2575 BUS[5].n16 BUS[5].t10 0.4555
R2576 BUS[5].n16 BUS[5].t18 0.4555
R2577 BUS[5].n14 BUS[5].t17 0.4555
R2578 BUS[5].n14 BUS[5].t8 0.4555
R2579 BUS[5].n12 BUS[5].t7 0.4555
R2580 BUS[5].n12 BUS[5].t15 0.4555
R2581 BUS[5].n10 BUS[5].t20 0.4555
R2582 BUS[5].n10 BUS[5].t22 0.4555
R2583 BUS[5].n8 BUS[5].t9 0.4555
R2584 BUS[5].n8 BUS[5].t12 0.4555
R2585 BUS[5].n7 BUS[5].t11 0.4555
R2586 BUS[5].n7 BUS[5].t19 0.4555
R2587 BUS[5].n5 BUS[5].t6 0.4555
R2588 BUS[5].n5 BUS[5].t14 0.4555
R2589 BUS[5].n0 BUS[5].t3 0.41
R2590 BUS[5].n0 BUS[5].t1 0.41
R2591 BUS[5].n1 BUS[5].t2 0.41
R2592 BUS[5].n1 BUS[5].t5 0.41
R2593 BUS[5].n3 BUS[5].t4 0.41
R2594 BUS[5].n3 BUS[5].t0 0.41
R2595 BUS[5].n4 BUS[5].n2 0.3605
R2596 BUS[5].n11 BUS[5].n9 0.3605
R2597 BUS[5].n13 BUS[5].n11 0.3605
R2598 BUS[5].n15 BUS[5].n13 0.3605
R2599 BUS[5].n17 BUS[5].n15 0.3605
R2600 BUS[5].n19 BUS[5].n17 0.3605
R2601 BUS[5].n21 BUS[5].n19 0.3605
R2602 BUS[5].n22 BUS[5].n6 0.203
R2603 BUS[5] BUS[5].n22 0.0430197
R2604 BUS[5].n22 BUS[5].n21 0.015125
R2605 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.7994
R2606 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R2607 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R2608 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R2609 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R2610 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R2611 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R2612 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R2613 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2614 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R2615 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R2616 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R2617 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R2618 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R2619 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R2620 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R2621 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R2622 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R2623 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R2624 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R2625 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R2626 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R2627 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R2628 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R2629 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R2630 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R2631 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R2632 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R2633 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R2634 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R2635 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R2636 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R2637 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R2638 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R2639 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R2640 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R2641 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R2642 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R2643 BUS[6].n2 BUS[6].n0 15.3751
R2644 BUS[6].n9 BUS[6].n7 15.2168
R2645 BUS[6].n2 BUS[6].n1 15.0151
R2646 BUS[6].n4 BUS[6].n3 15.0151
R2647 BUS[6].n21 BUS[6].n20 14.8568
R2648 BUS[6].n19 BUS[6].n18 14.8568
R2649 BUS[6].n17 BUS[6].n16 14.8568
R2650 BUS[6].n15 BUS[6].n14 14.8568
R2651 BUS[6].n13 BUS[6].n12 14.8568
R2652 BUS[6].n11 BUS[6].n10 14.8568
R2653 BUS[6].n9 BUS[6].n8 14.8568
R2654 BUS[6].n6 BUS[6].n5 14.8568
R2655 BUS[6].n22 BUS[6] 0.921051
R2656 BUS[6].n6 BUS[6].n4 0.8825
R2657 BUS[6].n20 BUS[6].t20 0.4555
R2658 BUS[6].n20 BUS[6].t11 0.4555
R2659 BUS[6].n18 BUS[6].t16 0.4555
R2660 BUS[6].n18 BUS[6].t23 0.4555
R2661 BUS[6].n16 BUS[6].t22 0.4555
R2662 BUS[6].n16 BUS[6].t13 0.4555
R2663 BUS[6].n14 BUS[6].t12 0.4555
R2664 BUS[6].n14 BUS[6].t15 0.4555
R2665 BUS[6].n12 BUS[6].t7 0.4555
R2666 BUS[6].n12 BUS[6].t9 0.4555
R2667 BUS[6].n10 BUS[6].t8 0.4555
R2668 BUS[6].n10 BUS[6].t18 0.4555
R2669 BUS[6].n8 BUS[6].t17 0.4555
R2670 BUS[6].n8 BUS[6].t6 0.4555
R2671 BUS[6].n7 BUS[6].t10 0.4555
R2672 BUS[6].n7 BUS[6].t14 0.4555
R2673 BUS[6].n5 BUS[6].t19 0.4555
R2674 BUS[6].n5 BUS[6].t21 0.4555
R2675 BUS[6].n0 BUS[6].t5 0.41
R2676 BUS[6].n0 BUS[6].t0 0.41
R2677 BUS[6].n1 BUS[6].t1 0.41
R2678 BUS[6].n1 BUS[6].t3 0.41
R2679 BUS[6].n3 BUS[6].t2 0.41
R2680 BUS[6].n3 BUS[6].t4 0.41
R2681 BUS[6].n4 BUS[6].n2 0.3605
R2682 BUS[6].n11 BUS[6].n9 0.3605
R2683 BUS[6].n13 BUS[6].n11 0.3605
R2684 BUS[6].n15 BUS[6].n13 0.3605
R2685 BUS[6].n17 BUS[6].n15 0.3605
R2686 BUS[6].n19 BUS[6].n17 0.3605
R2687 BUS[6].n21 BUS[6].n19 0.3605
R2688 BUS[6].n22 BUS[6].n6 0.203
R2689 BUS[6] BUS[6].n22 0.0430197
R2690 BUS[6].n22 BUS[6].n21 0.015125
R2691 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.7994
R2692 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R2693 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R2694 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R2695 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R2696 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R2697 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R2698 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R2699 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R2700 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R2701 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R2702 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R2703 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2704 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R2705 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R2706 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R2707 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R2708 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R2709 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R2710 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R2711 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R2712 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R2713 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R2714 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R2715 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R2716 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R2717 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R2718 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R2719 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R2720 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R2721 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R2722 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R2723 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R2724 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R2725 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R2726 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R2727 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R2728 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R2729 BUS[4].n2 BUS[4].n0 15.3751
R2730 BUS[4].n9 BUS[4].n7 15.2168
R2731 BUS[4].n2 BUS[4].n1 15.0151
R2732 BUS[4].n4 BUS[4].n3 15.0151
R2733 BUS[4].n21 BUS[4].n20 14.8568
R2734 BUS[4].n19 BUS[4].n18 14.8568
R2735 BUS[4].n17 BUS[4].n16 14.8568
R2736 BUS[4].n15 BUS[4].n14 14.8568
R2737 BUS[4].n13 BUS[4].n12 14.8568
R2738 BUS[4].n11 BUS[4].n10 14.8568
R2739 BUS[4].n9 BUS[4].n8 14.8568
R2740 BUS[4].n6 BUS[4].n5 14.8568
R2741 BUS[4].n22 BUS[4] 0.921051
R2742 BUS[4].n6 BUS[4].n4 0.8825
R2743 BUS[4].n20 BUS[4].t4 0.4555
R2744 BUS[4].n20 BUS[4].t12 0.4555
R2745 BUS[4].n18 BUS[4].t11 0.4555
R2746 BUS[4].n18 BUS[4].t2 0.4555
R2747 BUS[4].n16 BUS[4].t6 0.4555
R2748 BUS[4].n16 BUS[4].t3 0.4555
R2749 BUS[4].n14 BUS[4].t14 0.4555
R2750 BUS[4].n14 BUS[4].t17 0.4555
R2751 BUS[4].n12 BUS[4].t16 0.4555
R2752 BUS[4].n12 BUS[4].t5 0.4555
R2753 BUS[4].n10 BUS[4].t10 0.4555
R2754 BUS[4].n10 BUS[4].t13 0.4555
R2755 BUS[4].n8 BUS[4].t0 0.4555
R2756 BUS[4].n8 BUS[4].t8 0.4555
R2757 BUS[4].n7 BUS[4].t7 0.4555
R2758 BUS[4].n7 BUS[4].t9 0.4555
R2759 BUS[4].n5 BUS[4].t15 0.4555
R2760 BUS[4].n5 BUS[4].t1 0.4555
R2761 BUS[4].n0 BUS[4].t19 0.41
R2762 BUS[4].n0 BUS[4].t21 0.41
R2763 BUS[4].n1 BUS[4].t20 0.41
R2764 BUS[4].n1 BUS[4].t23 0.41
R2765 BUS[4].n3 BUS[4].t22 0.41
R2766 BUS[4].n3 BUS[4].t18 0.41
R2767 BUS[4].n4 BUS[4].n2 0.3605
R2768 BUS[4].n11 BUS[4].n9 0.3605
R2769 BUS[4].n13 BUS[4].n11 0.3605
R2770 BUS[4].n15 BUS[4].n13 0.3605
R2771 BUS[4].n17 BUS[4].n15 0.3605
R2772 BUS[4].n19 BUS[4].n17 0.3605
R2773 BUS[4].n21 BUS[4].n19 0.3605
R2774 BUS[4].n22 BUS[4].n6 0.203
R2775 BUS[4] BUS[4].n22 0.0430197
R2776 BUS[4].n22 BUS[4].n21 0.015125
R2777 PHI_2.n17 PHI_2.t19 26.4265
R2778 PHI_2.n15 PHI_2.t9 26.4265
R2779 PHI_2.n13 PHI_2.t8 26.4265
R2780 PHI_2.n11 PHI_2.t16 26.4265
R2781 PHI_2.n9 PHI_2.t12 26.4265
R2782 PHI_2.n7 PHI_2.t6 26.4265
R2783 PHI_2.n5 PHI_2.t0 26.4265
R2784 PHI_2.n3 PHI_2.t15 26.4265
R2785 PHI_2.n1 PHI_2.t4 26.4265
R2786 PHI_2.n0 PHI_2.t18 26.4265
R2787 PHI_2.n17 PHI_2.t2 11.7657
R2788 PHI_2.n15 PHI_2.t13 11.7657
R2789 PHI_2.n13 PHI_2.t10 11.7657
R2790 PHI_2.n11 PHI_2.t5 11.7657
R2791 PHI_2.n9 PHI_2.t14 11.7657
R2792 PHI_2.n7 PHI_2.t7 11.7657
R2793 PHI_2.n5 PHI_2.t3 11.7657
R2794 PHI_2.n3 PHI_2.t17 11.7657
R2795 PHI_2.n1 PHI_2.t11 11.7657
R2796 PHI_2.n0 PHI_2.t1 11.7657
R2797 PHI_2.n18 PHI_2 9.23499
R2798 PHI_2.n16 PHI_2 9.23499
R2799 PHI_2.n14 PHI_2 9.23499
R2800 PHI_2.n12 PHI_2 9.23499
R2801 PHI_2.n10 PHI_2 9.23499
R2802 PHI_2.n8 PHI_2 9.23499
R2803 PHI_2.n6 PHI_2 9.23499
R2804 PHI_2.n4 PHI_2 9.23499
R2805 PHI_2.n2 PHI_2 9.23499
R2806 PHI_2 PHI_2.n17 8.04257
R2807 PHI_2 PHI_2.n15 8.04257
R2808 PHI_2 PHI_2.n13 8.04257
R2809 PHI_2 PHI_2.n11 8.04257
R2810 PHI_2 PHI_2.n9 8.04257
R2811 PHI_2 PHI_2.n7 8.04257
R2812 PHI_2 PHI_2.n5 8.04257
R2813 PHI_2 PHI_2.n3 8.04257
R2814 PHI_2 PHI_2.n1 8.04257
R2815 PHI_2 PHI_2.n0 8.04257
R2816 PHI_2.n2 PHI_2 3.0407
R2817 PHI_2.n4 PHI_2 3.0407
R2818 PHI_2.n6 PHI_2 3.0407
R2819 PHI_2.n8 PHI_2 3.0407
R2820 PHI_2.n10 PHI_2 3.0407
R2821 PHI_2.n12 PHI_2 3.0407
R2822 PHI_2.n14 PHI_2 3.0407
R2823 PHI_2.n16 PHI_2 3.0407
R2824 PHI_2.n18 PHI_2 3.0407
R2825 PHI_2 PHI_2.n2 2.5763
R2826 PHI_2 PHI_2.n4 2.5763
R2827 PHI_2 PHI_2.n6 2.5763
R2828 PHI_2 PHI_2.n8 2.5763
R2829 PHI_2 PHI_2.n10 2.5763
R2830 PHI_2 PHI_2.n12 2.5763
R2831 PHI_2 PHI_2.n14 2.5763
R2832 PHI_2 PHI_2.n16 2.5763
R2833 PHI_2 PHI_2.n18 2.5763
R2834 BUS[8].n2 BUS[8].n0 15.3751
R2835 BUS[8].n9 BUS[8].n7 15.2168
R2836 BUS[8].n2 BUS[8].n1 15.0151
R2837 BUS[8].n4 BUS[8].n3 15.0151
R2838 BUS[8].n21 BUS[8].n20 14.8568
R2839 BUS[8].n19 BUS[8].n18 14.8568
R2840 BUS[8].n17 BUS[8].n16 14.8568
R2841 BUS[8].n15 BUS[8].n14 14.8568
R2842 BUS[8].n13 BUS[8].n12 14.8568
R2843 BUS[8].n11 BUS[8].n10 14.8568
R2844 BUS[8].n9 BUS[8].n8 14.8568
R2845 BUS[8].n6 BUS[8].n5 14.8568
R2846 BUS[8].n22 BUS[8] 0.921051
R2847 BUS[8].n6 BUS[8].n4 0.8825
R2848 BUS[8].n20 BUS[8].t4 0.4555
R2849 BUS[8].n20 BUS[8].t17 0.4555
R2850 BUS[8].n18 BUS[8].t18 0.4555
R2851 BUS[8].n18 BUS[8].t13 0.4555
R2852 BUS[8].n16 BUS[8].t21 0.4555
R2853 BUS[8].n16 BUS[8].t22 0.4555
R2854 BUS[8].n14 BUS[8].t15 0.4555
R2855 BUS[8].n14 BUS[8].t3 0.4555
R2856 BUS[8].n12 BUS[8].t11 0.4555
R2857 BUS[8].n12 BUS[8].t2 0.4555
R2858 BUS[8].n10 BUS[8].t19 0.4555
R2859 BUS[8].n10 BUS[8].t16 0.4555
R2860 BUS[8].n8 BUS[8].t0 0.4555
R2861 BUS[8].n8 BUS[8].t23 0.4555
R2862 BUS[8].n7 BUS[8].t20 0.4555
R2863 BUS[8].n7 BUS[8].t1 0.4555
R2864 BUS[8].n5 BUS[8].t12 0.4555
R2865 BUS[8].n5 BUS[8].t14 0.4555
R2866 BUS[8].n0 BUS[8].t5 0.41
R2867 BUS[8].n0 BUS[8].t9 0.41
R2868 BUS[8].n1 BUS[8].t8 0.41
R2869 BUS[8].n1 BUS[8].t10 0.41
R2870 BUS[8].n3 BUS[8].t6 0.41
R2871 BUS[8].n3 BUS[8].t7 0.41
R2872 BUS[8].n4 BUS[8].n2 0.3605
R2873 BUS[8].n11 BUS[8].n9 0.3605
R2874 BUS[8].n13 BUS[8].n11 0.3605
R2875 BUS[8].n15 BUS[8].n13 0.3605
R2876 BUS[8].n17 BUS[8].n15 0.3605
R2877 BUS[8].n19 BUS[8].n17 0.3605
R2878 BUS[8].n21 BUS[8].n19 0.3605
R2879 BUS[8].n22 BUS[8].n6 0.203
R2880 BUS[8] BUS[8].n22 0.0430197
R2881 BUS[8].n22 BUS[8].n21 0.015125
R2882 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.7994
R2883 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R2884 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R2885 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R2886 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R2887 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R2888 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R2889 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R2890 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R2891 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R2892 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R2893 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R2894 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R2895 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R2896 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R2897 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R2898 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R2899 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R2900 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R2901 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R2902 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R2903 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R2904 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R2905 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R2906 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R2907 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R2908 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R2909 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R2910 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R2911 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R2912 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R2913 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R2914 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R2915 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R2916 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R2917 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R2918 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R2919 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R2920 BUS[9].n2 BUS[9].n0 15.3751
R2921 BUS[9].n9 BUS[9].n7 15.2168
R2922 BUS[9].n2 BUS[9].n1 15.0151
R2923 BUS[9].n4 BUS[9].n3 15.0151
R2924 BUS[9].n21 BUS[9].n20 14.8568
R2925 BUS[9].n19 BUS[9].n18 14.8568
R2926 BUS[9].n17 BUS[9].n16 14.8568
R2927 BUS[9].n15 BUS[9].n14 14.8568
R2928 BUS[9].n13 BUS[9].n12 14.8568
R2929 BUS[9].n11 BUS[9].n10 14.8568
R2930 BUS[9].n9 BUS[9].n8 14.8568
R2931 BUS[9].n6 BUS[9].n5 14.8568
R2932 BUS[9].n22 BUS[9] 0.921051
R2933 BUS[9].n6 BUS[9].n4 0.8825
R2934 BUS[9].n20 BUS[9].t6 0.4555
R2935 BUS[9].n20 BUS[9].t17 0.4555
R2936 BUS[9].n18 BUS[9].t7 0.4555
R2937 BUS[9].n18 BUS[9].t22 0.4555
R2938 BUS[9].n16 BUS[9].t19 0.4555
R2939 BUS[9].n16 BUS[9].t20 0.4555
R2940 BUS[9].n14 BUS[9].t16 0.4555
R2941 BUS[9].n14 BUS[9].t2 0.4555
R2942 BUS[9].n12 BUS[9].t3 0.4555
R2943 BUS[9].n12 BUS[9].t4 0.4555
R2944 BUS[9].n10 BUS[9].t8 0.4555
R2945 BUS[9].n10 BUS[9].t23 0.4555
R2946 BUS[9].n8 BUS[9].t1 0.4555
R2947 BUS[9].n8 BUS[9].t21 0.4555
R2948 BUS[9].n7 BUS[9].t18 0.4555
R2949 BUS[9].n7 BUS[9].t0 0.4555
R2950 BUS[9].n5 BUS[9].t15 0.4555
R2951 BUS[9].n5 BUS[9].t5 0.4555
R2952 BUS[9].n0 BUS[9].t9 0.41
R2953 BUS[9].n0 BUS[9].t10 0.41
R2954 BUS[9].n1 BUS[9].t12 0.41
R2955 BUS[9].n1 BUS[9].t14 0.41
R2956 BUS[9].n3 BUS[9].t13 0.41
R2957 BUS[9].n3 BUS[9].t11 0.41
R2958 BUS[9].n4 BUS[9].n2 0.3605
R2959 BUS[9].n11 BUS[9].n9 0.3605
R2960 BUS[9].n13 BUS[9].n11 0.3605
R2961 BUS[9].n15 BUS[9].n13 0.3605
R2962 BUS[9].n17 BUS[9].n15 0.3605
R2963 BUS[9].n19 BUS[9].n17 0.3605
R2964 BUS[9].n21 BUS[9].n19 0.3605
R2965 BUS[9].n22 BUS[9].n6 0.203
R2966 BUS[9] BUS[9].n22 0.0430197
R2967 BUS[9].n22 BUS[9].n21 0.015125
R2968 enable.n18 enable.t10 19.9538
R2969 enable.n16 enable.t11 19.9538
R2970 enable.n14 enable.t4 19.9538
R2971 enable.n12 enable.t8 19.9538
R2972 enable.n10 enable.t17 19.9538
R2973 enable.n8 enable.t19 19.9538
R2974 enable.n6 enable.t5 19.9538
R2975 enable.n4 enable.t15 19.9538
R2976 enable.n2 enable.t0 19.9538
R2977 enable.n0 enable.t7 19.9538
R2978 enable.n18 enable.t2 17.3015
R2979 enable.n16 enable.t3 17.3015
R2980 enable.n14 enable.t14 17.3015
R2981 enable.n12 enable.t18 17.3015
R2982 enable.n10 enable.t6 17.3015
R2983 enable.n8 enable.t12 17.3015
R2984 enable.n6 enable.t16 17.3015
R2985 enable.n4 enable.t9 17.3015
R2986 enable.n2 enable.t13 17.3015
R2987 enable.n0 enable.t1 17.3015
R2988 enable enable.n19 10.8498
R2989 enable.n19 enable.n18 8.0005
R2990 enable.n17 enable.n16 8.0005
R2991 enable.n15 enable.n14 8.0005
R2992 enable.n13 enable.n12 8.0005
R2993 enable.n11 enable.n10 8.0005
R2994 enable.n9 enable.n8 8.0005
R2995 enable.n7 enable.n6 8.0005
R2996 enable.n5 enable.n4 8.0005
R2997 enable.n3 enable.n2 8.0005
R2998 enable.n1 enable.n0 8.0005
R2999 enable enable.n20 6.01421
R3000 enable enable.n21 6.01421
R3001 enable enable.n22 6.01421
R3002 enable enable.n23 6.01421
R3003 enable enable.n24 6.01421
R3004 enable enable.n25 6.01421
R3005 enable enable.n26 6.01421
R3006 enable enable.n27 6.01421
R3007 enable enable.n28 6.01421
R3008 enable.n20 enable.n17 4.8361
R3009 enable.n21 enable.n15 4.8361
R3010 enable.n22 enable.n13 4.8361
R3011 enable.n23 enable.n11 4.8361
R3012 enable.n24 enable.n9 4.8361
R3013 enable.n25 enable.n7 4.8361
R3014 enable.n26 enable.n5 4.8361
R3015 enable.n27 enable.n3 4.8361
R3016 enable.n28 enable.n1 4.8361
R3017 enable.n20 enable 1.07965
R3018 enable.n21 enable 1.07965
R3019 enable.n22 enable 1.07965
R3020 enable.n23 enable 1.07965
R3021 enable.n24 enable 1.07965
R3022 enable.n25 enable 1.07965
R3023 enable.n26 enable 1.07965
R3024 enable.n27 enable 1.07965
R3025 enable.n28 enable 1.07965
R3026 enable.n19 enable 0.00742308
R3027 enable.n17 enable 0.00742308
R3028 enable.n15 enable 0.00742308
R3029 enable.n13 enable 0.00742308
R3030 enable.n11 enable 0.00742308
R3031 enable.n9 enable 0.00742308
R3032 enable.n7 enable 0.00742308
R3033 enable.n5 enable 0.00742308
R3034 enable.n3 enable 0.00742308
R3035 enable.n1 enable 0.00742308
R3036 PHI_1.n17 PHI_1.t2 26.4265
R3037 PHI_1.n15 PHI_1.t9 26.4265
R3038 PHI_1.n13 PHI_1.t1 26.4265
R3039 PHI_1.n11 PHI_1.t12 26.4265
R3040 PHI_1.n9 PHI_1.t11 26.4265
R3041 PHI_1.n7 PHI_1.t19 26.4265
R3042 PHI_1.n5 PHI_1.t16 26.4265
R3043 PHI_1.n3 PHI_1.t8 26.4265
R3044 PHI_1.n1 PHI_1.t4 26.4265
R3045 PHI_1.n0 PHI_1.t18 26.4265
R3046 PHI_1.n17 PHI_1.t3 11.7657
R3047 PHI_1.n15 PHI_1.t13 11.7657
R3048 PHI_1.n13 PHI_1.t5 11.7657
R3049 PHI_1.n11 PHI_1.t15 11.7657
R3050 PHI_1.n9 PHI_1.t14 11.7657
R3051 PHI_1.n7 PHI_1.t7 11.7657
R3052 PHI_1.n5 PHI_1.t17 11.7657
R3053 PHI_1.n3 PHI_1.t10 11.7657
R3054 PHI_1.n1 PHI_1.t6 11.7657
R3055 PHI_1.n0 PHI_1.t0 11.7657
R3056 PHI_1.n18 PHI_1 9.56151
R3057 PHI_1.n16 PHI_1 9.56151
R3058 PHI_1.n14 PHI_1 9.56151
R3059 PHI_1.n12 PHI_1 9.56151
R3060 PHI_1.n10 PHI_1 9.56151
R3061 PHI_1.n8 PHI_1 9.56151
R3062 PHI_1.n6 PHI_1 9.56151
R3063 PHI_1.n4 PHI_1 9.56151
R3064 PHI_1.n2 PHI_1 9.56151
R3065 PHI_1 PHI_1.n17 8.04713
R3066 PHI_1 PHI_1.n15 8.04713
R3067 PHI_1 PHI_1.n13 8.04713
R3068 PHI_1 PHI_1.n11 8.04713
R3069 PHI_1 PHI_1.n9 8.04713
R3070 PHI_1 PHI_1.n7 8.04713
R3071 PHI_1 PHI_1.n5 8.04713
R3072 PHI_1 PHI_1.n3 8.04713
R3073 PHI_1 PHI_1.n1 8.04713
R3074 PHI_1 PHI_1.n0 8.04713
R3075 PHI_1.n2 PHI_1 5.2583
R3076 PHI_1.n4 PHI_1 5.2583
R3077 PHI_1.n6 PHI_1 5.2583
R3078 PHI_1.n8 PHI_1 5.2583
R3079 PHI_1.n10 PHI_1 5.2583
R3080 PHI_1.n12 PHI_1 5.2583
R3081 PHI_1.n14 PHI_1 5.2583
R3082 PHI_1.n16 PHI_1 5.2583
R3083 PHI_1.n18 PHI_1 5.2583
R3084 PHI_1 PHI_1.n2 0.3587
R3085 PHI_1 PHI_1.n4 0.3587
R3086 PHI_1 PHI_1.n6 0.3587
R3087 PHI_1 PHI_1.n8 0.3587
R3088 PHI_1 PHI_1.n10 0.3587
R3089 PHI_1 PHI_1.n12 0.3587
R3090 PHI_1 PHI_1.n14 0.3587
R3091 PHI_1 PHI_1.n16 0.3587
R3092 PHI_1 PHI_1.n18 0.3587
R3093 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.7994
R3094 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R3095 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R3096 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R3097 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R3098 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R3099 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R3100 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R3101 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R3102 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R3103 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R3104 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R3105 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R3106 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R3107 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R3108 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R3109 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R3110 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R3111 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R3112 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R3113 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R3114 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R3115 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R3116 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R3117 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R3118 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R3119 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R3120 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R3121 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R3122 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R3123 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R3124 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R3125 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R3126 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R3127 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R3128 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R3129 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R3130 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R3131 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.7994
R3132 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R3133 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R3134 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R3135 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R3136 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R3137 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R3138 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R3139 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R3140 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R3141 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R3142 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R3143 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R3144 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R3145 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R3146 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R3147 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R3148 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R3149 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R3150 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R3151 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R3152 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R3153 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R3154 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R3155 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R3156 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R3157 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R3158 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R3159 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R3160 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R3161 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R3162 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R3163 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R3164 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R3165 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R3166 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R3167 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R3168 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R3169 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.7994
R3170 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R3171 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R3172 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R3173 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R3174 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R3175 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R3176 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R3177 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R3178 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R3179 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R3180 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R3181 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R3182 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R3183 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.6148
R3184 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R3185 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R3186 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R3187 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R3188 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R3189 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R3190 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R3191 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R3192 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R3193 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R3194 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R3195 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R3196 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R3197 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R3198 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R3199 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R3200 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R3201 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R3202 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R3203 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R3204 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R3205 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R3206 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R3207 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 71.7994
R3208 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 71.6148
R3209 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 71.6148
R3210 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 71.6148
R3211 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 71.6148
R3212 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 71.6148
R3213 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 71.6148
R3214 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 71.6148
R3215 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 71.6148
R3216 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 71.6148
R3217 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 71.6148
R3218 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 71.6148
R3219 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 71.6148
R3220 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 71.6148
R3221 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 71.6148
R3222 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 71.6148
R3223 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 71.6148
R3224 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 71.6148
R3225 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 11.4757
R3226 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 4.63372
R3227 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 3.85252
R3228 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 0.402556
R3229 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 0.185115
R3230 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 0.185115
R3231 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 0.185115
R3232 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 0.185115
R3233 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 0.185115
R3234 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 0.185115
R3235 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 0.185115
R3236 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 0.185115
R3237 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 0.185115
R3238 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 0.185115
R3239 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 0.185115
R3240 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 0.185115
R3241 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 0.185115
R3242 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 0.185115
R3243 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 0.185115
R3244 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 0.185115
R3245 BUS[3].n2 BUS[3].n0 15.3751
R3246 BUS[3].n9 BUS[3].n7 15.2168
R3247 BUS[3].n2 BUS[3].n1 15.0151
R3248 BUS[3].n4 BUS[3].n3 15.0151
R3249 BUS[3].n21 BUS[3].n20 14.8568
R3250 BUS[3].n19 BUS[3].n18 14.8568
R3251 BUS[3].n17 BUS[3].n16 14.8568
R3252 BUS[3].n15 BUS[3].n14 14.8568
R3253 BUS[3].n13 BUS[3].n12 14.8568
R3254 BUS[3].n11 BUS[3].n10 14.8568
R3255 BUS[3].n9 BUS[3].n8 14.8568
R3256 BUS[3].n6 BUS[3].n5 14.8568
R3257 BUS[3].n22 BUS[3] 0.921051
R3258 BUS[3].n6 BUS[3].n4 0.8825
R3259 BUS[3].n20 BUS[3].t16 0.4555
R3260 BUS[3].n20 BUS[3].t1 0.4555
R3261 BUS[3].n18 BUS[3].t0 0.4555
R3262 BUS[3].n18 BUS[3].t10 0.4555
R3263 BUS[3].n16 BUS[3].t9 0.4555
R3264 BUS[3].n16 BUS[3].t15 0.4555
R3265 BUS[3].n14 BUS[3].t3 0.4555
R3266 BUS[3].n14 BUS[3].t6 0.4555
R3267 BUS[3].n12 BUS[3].t12 0.4555
R3268 BUS[3].n12 BUS[3].t13 0.4555
R3269 BUS[3].n10 BUS[3].t17 0.4555
R3270 BUS[3].n10 BUS[3].t2 0.4555
R3271 BUS[3].n8 BUS[3].t7 0.4555
R3272 BUS[3].n8 BUS[3].t11 0.4555
R3273 BUS[3].n7 BUS[3].t14 0.4555
R3274 BUS[3].n7 BUS[3].t4 0.4555
R3275 BUS[3].n5 BUS[3].t5 0.4555
R3276 BUS[3].n5 BUS[3].t8 0.4555
R3277 BUS[3].n0 BUS[3].t19 0.41
R3278 BUS[3].n0 BUS[3].t22 0.41
R3279 BUS[3].n1 BUS[3].t21 0.41
R3280 BUS[3].n1 BUS[3].t23 0.41
R3281 BUS[3].n3 BUS[3].t20 0.41
R3282 BUS[3].n3 BUS[3].t18 0.41
R3283 BUS[3].n4 BUS[3].n2 0.3605
R3284 BUS[3].n11 BUS[3].n9 0.3605
R3285 BUS[3].n13 BUS[3].n11 0.3605
R3286 BUS[3].n15 BUS[3].n13 0.3605
R3287 BUS[3].n17 BUS[3].n15 0.3605
R3288 BUS[3].n19 BUS[3].n17 0.3605
R3289 BUS[3].n21 BUS[3].n19 0.3605
R3290 BUS[3].n22 BUS[3].n6 0.203
R3291 BUS[3] BUS[3].n22 0.0430197
R3292 BUS[3].n22 BUS[3].n21 0.015125
R3293 BUS[10].n2 BUS[10].n0 15.3751
R3294 BUS[10].n9 BUS[10].n7 15.2168
R3295 BUS[10].n2 BUS[10].n1 15.0151
R3296 BUS[10].n4 BUS[10].n3 15.0151
R3297 BUS[10].n21 BUS[10].n20 14.8568
R3298 BUS[10].n19 BUS[10].n18 14.8568
R3299 BUS[10].n17 BUS[10].n16 14.8568
R3300 BUS[10].n15 BUS[10].n14 14.8568
R3301 BUS[10].n13 BUS[10].n12 14.8568
R3302 BUS[10].n11 BUS[10].n10 14.8568
R3303 BUS[10].n9 BUS[10].n8 14.8568
R3304 BUS[10].n6 BUS[10].n5 14.8568
R3305 BUS[10].n22 BUS[10] 0.921051
R3306 BUS[10].n6 BUS[10].n4 0.8825
R3307 BUS[10].n20 BUS[10].t16 0.4555
R3308 BUS[10].n20 BUS[10].t20 0.4555
R3309 BUS[10].n18 BUS[10].t10 0.4555
R3310 BUS[10].n18 BUS[10].t13 0.4555
R3311 BUS[10].n16 BUS[10].t12 0.4555
R3312 BUS[10].n16 BUS[10].t22 0.4555
R3313 BUS[10].n14 BUS[10].t21 0.4555
R3314 BUS[10].n14 BUS[10].t9 0.4555
R3315 BUS[10].n12 BUS[10].t7 0.4555
R3316 BUS[10].n12 BUS[10].t18 0.4555
R3317 BUS[10].n10 BUS[10].t15 0.4555
R3318 BUS[10].n10 BUS[10].t19 0.4555
R3319 BUS[10].n8 BUS[10].t23 0.4555
R3320 BUS[10].n8 BUS[10].t6 0.4555
R3321 BUS[10].n7 BUS[10].t11 0.4555
R3322 BUS[10].n7 BUS[10].t14 0.4555
R3323 BUS[10].n5 BUS[10].t8 0.4555
R3324 BUS[10].n5 BUS[10].t17 0.4555
R3325 BUS[10].n0 BUS[10].t3 0.41
R3326 BUS[10].n0 BUS[10].t4 0.41
R3327 BUS[10].n1 BUS[10].t5 0.41
R3328 BUS[10].n1 BUS[10].t1 0.41
R3329 BUS[10].n3 BUS[10].t0 0.41
R3330 BUS[10].n3 BUS[10].t2 0.41
R3331 BUS[10].n4 BUS[10].n2 0.3605
R3332 BUS[10].n11 BUS[10].n9 0.3605
R3333 BUS[10].n13 BUS[10].n11 0.3605
R3334 BUS[10].n15 BUS[10].n13 0.3605
R3335 BUS[10].n17 BUS[10].n15 0.3605
R3336 BUS[10].n19 BUS[10].n17 0.3605
R3337 BUS[10].n21 BUS[10].n19 0.3605
R3338 BUS[10].n22 BUS[10].n6 0.203
R3339 BUS[10] BUS[10].n22 0.0430197
R3340 BUS[10].n22 BUS[10].n21 0.015125
R3341 d_out.n0 d_out.t2 21.1948
R3342 d_out.n0 d_out.t3 16.0605
R3343 d_out d_out.n3 9.16609
R3344 d_out.n2 d_out.n1 9.0005
R3345 d_out.n1 d_out.n0 8.12012
R3346 d_out.n2 d_out 5.47636
R3347 d_out.n3 d_out.t0 4.5901
R3348 d_out d_out.t1 3.91488
R3349 d_out.n3 d_out 0.150731
R3350 d_out d_out.n2 0.13775
R3351 d_out.n1 d_out 0.00840541
R3352 D_in.n0 D_in.t0 29.4195
R3353 D_in.n0 D_in.t1 11.4372
R3354 D_in D_in.n1 9.95
R3355 D_in.n1 D_in.n0 8.0005
R3356 D_in.n1 D_in 0.102506
C0 a_47136_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1 a_41140_1577# enable 0.00579f
C2 a_33672_1562# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C3 a_18728_1562# a_19196_1580# 0.30528f
C4 swmatrix_Tgate_8.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C5 a_28416_2122# vdd 0.55944f
C6 a_25952_2122# vdd 0.56482f
C7 ShiftReg_row_10_2$1_0.Q[7] a_44156_1580# 0.36203f
C8 a_15936_2122# a_16280_2002# 0.57845f
C9 swmatrix_Tgate_4.gated_control enable 0.50846f
C10 a_47380_1577# pin 0
C11 a_14952_1562# a_15420_1580# 0.30528f
C12 a_13472_2122# a_12956_1580# 0.30053f
C13 a_26296_2002# swmatrix_Tgate_5.gated_control 0.01121f
C14 swmatrix_Tgate_7.gated_control pin 1.23291f
C15 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_8.gated_control 0.17277f
C16 a_47480_2002# vdd 0.32887f
C17 a_44156_1580# vdd 0.42253f
C18 a_59616_2122# PHI_2 0.04011f
C19 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_53720_2002# 0.00242f
C20 a_15420_1580# pin 0.00113f
C21 a_57152_2122# PHI_2 0.04895f
C22 a_50396_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C23 a_28620_2122# BUS[5] 0.00104f
C24 a_14952_1562# pin 0.00138f
C25 a_9696_2122# BUS[2] 0.01571f
C26 a_25804_2122# BUS[5] 0
C27 a_7232_2122# BUS[2] 0.0191f
C28 a_28268_2122# enable 0.00101f
C29 a_54841_1539# BUS[9] 0
C30 a_1236_1577# BUS[1] 0
C31 a_2940_1580# PHI_2 0.07395f
C32 a_26296_2002# enable 0.05124f
C33 a_3660_2122# swmatrix_Tgate_9.gated_control 0
C34 a_59468_1577# enable 0.0022f
C35 a_35000_2002# a_34860_2122# 0.00109f
C36 a_32192_2122# a_32044_1577# 0
C37 a_9940_1577# BUS[2] 0
C38 a_24968_1562# swmatrix_Tgate_7.gated_control 0.00493f
C39 a_31676_1580# a_32044_2122# 0.00294f
C40 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C41 a_32536_2002# pin 0.00146f
C42 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_3.gated_control 0.22418f
C43 a_44916_1577# enable 0.00577f
C44 a_34656_2122# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C45 a_32192_2122# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C46 a_18728_1562# a_21192_1562# 0
C47 a_44876_2122# enable 0.00368f
C48 ShiftReg_row_10_2$1_0.Q[2] vdd 0.57779f
C49 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C50 a_51156_1577# pin 0
C51 a_40380_1580# a_40748_1577# 0.00194f
C52 a_18728_1562# enable 0.08752f
C53 swmatrix_Tgate_3.gated_control BUS[8] 0.86843f
C54 a_15936_2122# a_15420_1580# 0.30053f
C55 a_41240_2002# a_41140_1577# 0
C56 a_14952_1562# a_15936_2122# 0.07055f
C57 swmatrix_Tgate_1.gated_control vdd 1.84761f
C58 a_13472_2122# a_14952_1562# 0.00268f
C59 a_28760_2002# swmatrix_Tgate_5.gated_control 0.01014f
C60 a_25436_1580# swmatrix_Tgate_5.gated_control 0.00804f
C61 a_24968_1562# pin 0
C62 a_46620_1580# vdd 0.42496f
C63 a_46152_1562# vdd 1.0427f
C64 ShiftReg_row_10_2$1_0.Q[1] PHI_2 0.63578f
C65 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_52860_1580# 0.36162f
C66 a_52392_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C67 a_15936_2122# pin 0.00251f
C68 a_28268_2122# BUS[5] 0
C69 a_13472_2122# pin 0.00138f
C70 a_19916_2122# PHI_1 0.00534f
C71 a_26296_2002# BUS[5] 0.0117f
C72 a_53228_1577# BUS[9] 0
C73 a_28760_2002# enable 0.0522f
C74 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C75 a_3456_2122# PHI_2 0.04011f
C76 a_25436_1580# enable 0.05108f
C77 a_59860_1577# enable 0.00579f
C78 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[3] 0.10774f
C79 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_9.gated_control 0.33472f
C80 ShiftReg_row_10_2$1_0.Q[7] PHI_1 0.05798f
C81 a_32192_2122# a_32436_1577# 0.01595f
C82 a_35000_2002# pin 0
C83 a_31676_1580# a_32536_2002# 0.00888f
C84 a_31676_1580# pin 0
C85 a_32192_2122# a_32396_2122# 0.01151f
C86 ShiftReg_row_10_2$1_0.Q[8] a_49928_1562# 0.16779f
C87 a_44524_1577# swmatrix_Tgate_3.gated_control 0
C88 a_47340_2122# enable 0.00368f
C89 a_18728_1562# a_19712_2122# 0.07055f
C90 a_44524_2122# enable 0.00101f
C91 a_992_2122# vdd 0.56615f
C92 vdd PHI_1 9.89729f
C93 swmatrix_Tgate_5.gated_control swmatrix_Tgate_6.gated_control 0.01259f
C94 a_476_1580# PHI_1 0.0533f
C95 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C96 a_8_1562# a_1336_2002# 0.02403f
C97 a_992_2122# a_476_1580# 0.30053f
C98 ShiftReg_row_10_2$1_0.Q[7] a_44672_2122# 0.01552f
C99 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C100 pin BUS[1] 11.0721f
C101 a_40896_2122# a_40748_1577# 0
C102 a_56168_1562# vdd 1.00067f
C103 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C104 a_27900_1580# swmatrix_Tgate_5.gated_control 0.00668f
C105 swmatrix_Tgate_1.gated_control a_54841_1539# 0.00113f
C106 a_56168_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C107 a_27432_1562# swmatrix_Tgate_5.gated_control 0.00985f
C108 a_47136_2122# vdd 0.55944f
C109 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_3308_1577# 0
C110 a_44672_2122# vdd 0.56482f
C111 a_53720_2002# ShiftReg_row_10_2$1_0.Q[9] 0.25874f
C112 swmatrix_Tgate_2.gated_control PHI_2 0.31095f
C113 ShiftReg_row_10_2$1_0.Q[4] ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C114 a_22380_2122# PHI_1 0.00477f
C115 swmatrix_Tgate_6.gated_control enable 0.50846f
C116 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_53376_2122# 0.01536f
C117 a_19564_2122# PHI_1 0.00201f
C118 a_50912_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C119 a_28760_2002# BUS[5] 0.01161f
C120 a_12488_1562# swmatrix_Tgate_8.gated_control 0.00493f
C121 a_25436_1580# BUS[5] 0.00688f
C122 swmatrix_Tgate_8.gated_control PHI_2 0.31095f
C123 PHI_1 BUS[4] 0.09486f
C124 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C125 a_27432_1562# enable 0.08694f
C126 swmatrix_Tgate_0.gated_control pin 1.23291f
C127 ShiftReg_row_10_2$1_0.Q[3] ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C128 a_53620_1577# BUS[9] 0
C129 a_27900_1580# enable 0.05124f
C130 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_15788_1577# 0
C131 a_34140_1580# a_34508_2122# 0.00294f
C132 a_34656_2122# a_34860_2122# 0.01151f
C133 swmatrix_Tgate_2.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C134 a_3800_2002# swmatrix_Tgate_9.gated_control 0.01014f
C135 a_34140_1580# pin 0.00113f
C136 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_6248_1562# 0
C137 a_33672_1562# a_32536_2002# 0
C138 a_33672_1562# pin 0.00138f
C139 a_32192_2122# a_32044_2122# 0
C140 a_44916_1577# swmatrix_Tgate_3.gated_control 0
C141 a_46988_2122# enable 0.00101f
C142 a_44876_2122# swmatrix_Tgate_3.gated_control 0
C143 a_7436_2122# vdd 0.01506f
C144 a_45016_2002# enable 0.05124f
C145 a_40896_2122# a_41140_1577# 0.01595f
C146 a_2472_1562# PHI_1 0.01733f
C147 a_31208_1562# swmatrix_Tgate_6.gated_control 0.01486f
C148 a_992_2122# a_2472_1562# 0.00268f
C149 enable BUS[9] 0.2115f
C150 a_51256_2002# pin 0.00146f
C151 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C152 swmatrix_Tgate_1.gated_control a_53228_1577# 0
C153 a_28416_2122# swmatrix_Tgate_5.gated_control 0.01553f
C154 a_25952_2122# swmatrix_Tgate_5.gated_control 0.01496f
C155 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C156 swmatrix_Tgate_6.gated_control BUS[5] 0.00566f
C157 a_844_2122# vdd 0.00491f
C158 a_476_1580# a_844_2122# 0.00294f
C159 a_992_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C160 a_52860_1580# ShiftReg_row_10_2$1_0.Q[9] 0.00101f
C161 a_3800_2002# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00186f
C162 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C163 a_51256_2002# a_51156_1577# 0
C164 a_52392_1562# ShiftReg_row_10_2$1_0.Q[9] 0.00225f
C165 a_50396_1580# a_50764_1577# 0.00194f
C166 a_22028_2122# PHI_1 0.00164f
C167 a_51256_2002# a_51116_2122# 0.00109f
C168 a_37448_1562# enable 0.08752f
C169 a_27900_1580# BUS[5] 0.01336f
C170 a_20056_2002# PHI_1 0.01314f
C171 vdd BUS[10] 0.56053f
C172 a_27432_1562# BUS[5] 0.02637f
C173 a_12488_1562# PHI_2 0.02762f
C174 a_43688_1562# pin 0
C175 swmatrix_Tgate_3.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C176 a_4921_1539# enable 0.00398f
C177 a_28416_2122# enable 0.11443f
C178 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[10] 0.10774f
C179 ShiftReg_row_10_2$1_0.Q[3] a_17401_1539# 0.00241f
C180 a_37448_1562# a_38776_2002# 0.02403f
C181 a_25952_2122# enable 0.11055f
C182 swmatrix_Tgate_6.gated_control a_37916_1580# 0
C183 a_2940_1580# swmatrix_Tgate_9.gated_control 0.00668f
C184 ShiftReg_row_10_2$1_0.Q[3] BUS[3] 0.01695f
C185 a_34656_2122# a_34508_2122# 0
C186 a_34140_1580# a_35000_2002# 0.00888f
C187 a_33672_1562# a_35000_2002# 0.02403f
C188 a_34656_2122# pin 0.00251f
C189 a_32192_2122# a_32536_2002# 0.57845f
C190 a_33672_1562# a_31676_1580# 0
C191 PHI_2 BUS[7] 0.11252f
C192 a_32192_2122# pin 0.00138f
C193 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_29881_1539# 0.0097f
C194 a_38636_2122# PHI_1 0.00534f
C195 a_47340_2122# swmatrix_Tgate_3.gated_control 0
C196 a_47480_2002# enable 0.0522f
C197 a_44156_1580# enable 0.05108f
C198 a_9900_2122# vdd 0.01506f
C199 a_7084_2122# vdd 0.00491f
C200 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C201 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C202 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.01636f
C203 a_53720_2002# pin 0
C204 a_50396_1580# pin 0
C205 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C206 ShiftReg_row_10_2$1_0.Q[2] ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C207 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C208 swmatrix_Tgate_1.gated_control a_57004_1577# 0
C209 swmatrix_Tgate_1.gated_control a_53620_1577# 0
C210 a_23641_1539# PHI_2 0
C211 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C212 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C213 a_1336_2002# vdd 0.32604f
C214 a_1196_2122# PHI_1 0.00534f
C215 a_53376_2122# ShiftReg_row_10_2$1_0.Q[9] 0.11433f
C216 a_2940_1580# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00199f
C217 a_992_2122# a_1196_2122# 0.01151f
C218 a_476_1580# a_1336_2002# 0.00888f
C219 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_9.gated_control 0.22418f
C220 a_22520_2002# PHI_1 0.01261f
C221 a_19196_1580# PHI_1 0.0533f
C222 a_28416_2122# BUS[5] 0.01571f
C223 ShiftReg_row_10_2$1_0.Q[2] enable 0.513f
C224 a_25952_2122# BUS[5] 0.0191f
C225 a_37448_1562# a_37916_1580# 0.30528f
C226 a_3308_1577# enable 0.0022f
C227 a_3456_2122# swmatrix_Tgate_9.gated_control 0.01553f
C228 a_13324_1577# BUS[3] 0
C229 a_34656_2122# a_35000_2002# 0.57845f
C230 swmatrix_Tgate_1.gated_control enable 0.50846f
C231 a_24968_1562# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C232 a_41100_2122# PHI_1 0.00477f
C233 a_33672_1562# a_34140_1580# 0.30528f
C234 a_32192_2122# a_31676_1580# 0.30053f
C235 a_38284_2122# PHI_1 0.00201f
C236 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[5] 0.01102f
C237 a_46620_1580# enable 0.05124f
C238 a_45016_2002# swmatrix_Tgate_3.gated_control 0.01121f
C239 a_9548_2122# vdd 0.00491f
C240 a_46152_1562# enable 0.08694f
C241 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C242 a_7576_2002# vdd 0.32603f
C243 a_38284_1577# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C244 a_6248_1562# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C245 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00368f
C246 a_52860_1580# pin 0.00113f
C247 a_59100_1580# a_59468_1577# 0.00194f
C248 a_59960_2002# a_59860_1577# 0
C249 a_52392_1562# pin 0.00138f
C250 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C251 ShiftReg_row_10_2$1_0.Q[5] PHI_2 0.63578f
C252 a_22028_1577# PHI_2 0
C253 swmatrix_Tgate_5.gated_control PHI_1 0.01086f
C254 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C255 a_3456_2122# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00396f
C256 a_53720_2002# a_53580_2122# 0.00109f
C257 a_2472_1562# a_1336_2002# 0
C258 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C259 ShiftReg_row_10_2$1_0.Q[1] a_6248_1562# 0.16779f
C260 a_43688_1562# swmatrix_Tgate_0.gated_control 0.00493f
C261 a_50912_2122# a_50764_1577# 0
C262 a_21660_1580# PHI_1 0.01277f
C263 a_50396_1580# a_50764_2122# 0.00294f
C264 a_21192_1562# PHI_1 0.01733f
C265 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C266 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[4] 0
C267 a_7084_1577# enable 0.0022f
C268 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[10] 0
C269 ShiftReg_row_10_2$1_0.Q[3] a_19564_1577# 0
C270 a_3700_1577# enable 0.00579f
C271 swmatrix_Tgate_9.gated_control swmatrix_Tgate_8.gated_control 0.01259f
C272 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C273 a_992_2122# enable 0.11055f
C274 D_in PHI_2 0.34149f
C275 a_37448_1562# a_39912_1562# 0
C276 PHI_1 enable 0.59089f
C277 a_1336_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C278 a_13716_1577# BUS[3] 0
C279 a_34656_2122# a_34140_1580# 0.30053f
C280 a_13676_2122# BUS[3] 0
C281 a_40748_2122# PHI_1 0.00164f
C282 a_56168_1562# enable 0.08752f
C283 a_38776_2002# PHI_1 0.01314f
C284 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C285 a_33672_1562# a_34656_2122# 0.07055f
C286 a_32192_2122# a_33672_1562# 0.00268f
C287 a_47480_2002# swmatrix_Tgate_3.gated_control 0.01014f
C288 a_47136_2122# enable 0.11443f
C289 a_44156_1580# swmatrix_Tgate_3.gated_control 0.00804f
C290 a_10040_2002# vdd 0.32887f
C291 a_6716_1580# vdd 0.42253f
C292 a_44672_2122# enable 0.11055f
C293 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_4.gated_control 0.33472f
C294 a_53376_2122# pin 0.00251f
C295 a_38676_1577# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C296 a_49928_1562# BUS[9] 0.0057f
C297 pin BUS[2] 11.0719f
C298 a_59616_2122# a_59468_1577# 0
C299 a_57356_2122# PHI_1 0.00534f
C300 a_50912_2122# pin 0.00138f
C301 swmatrix_Tgate_4.gated_control swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C302 a_25804_1577# PHI_2 0
C303 swmatrix_Tgate_8.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00338f
C304 a_22420_1577# PHI_2 0
C305 a_31208_1562# PHI_1 0.70141f
C306 a_22176_2122# PHI_1 0.01804f
C307 a_50912_2122# a_51156_1577# 0.01595f
C308 a_19712_2122# PHI_1 0.01882f
C309 a_50912_2122# a_51116_2122# 0.01151f
C310 a_50396_1580# a_51256_2002# 0.00888f
C311 PHI_1 BUS[5] 0.09486f
C312 a_57004_1577# BUS[10] 0
C313 a_7476_1577# enable 0.00577f
C314 a_37448_1562# a_38432_2122# 0.07055f
C315 a_42361_1539# PHI_2 0
C316 a_6248_1562# swmatrix_Tgate_8.gated_control 0.01486f
C317 a_7436_2122# enable 0.00368f
C318 swmatrix_Tgate_9.gated_control PHI_2 0.31101f
C319 a_1336_2002# a_1196_2122# 0.00109f
C320 swmatrix_Tgate_3.gated_control swmatrix_Tgate_1.gated_control 0.01259f
C321 a_16140_2122# BUS[3] 0.00104f
C322 a_41240_2002# PHI_1 0.01261f
C323 a_13324_2122# BUS[3] 0
C324 a_37916_1580# PHI_1 0.0533f
C325 a_42361_1539# BUS[7] 0
C326 a_46620_1580# swmatrix_Tgate_3.gated_control 0.00668f
C327 a_46152_1562# swmatrix_Tgate_3.gated_control 0.00985f
C328 a_9180_1580# vdd 0.42496f
C329 a_844_2122# enable 0.00101f
C330 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_18728_1562# 0
C331 a_8712_1562# vdd 1.0427f
C332 swmatrix_Tgate_2.gated_control a_61081_1539# 0.00113f
C333 ShiftReg_row_10_2$1_0.Q[7] ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C334 enable BUS[10] 0.2115f
C335 a_59820_2122# PHI_1 0.00477f
C336 a_59616_2122# a_59860_1577# 0.01595f
C337 a_57004_2122# PHI_1 0.00201f
C338 ShiftReg_row_10_2$1_0.Q[3] vdd 0.57779f
C339 ShiftReg_row_10_2$1_0.Q[6] ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C340 a_26196_1577# PHI_2 0
C341 a_26156_2122# PHI_2 0.00411f
C342 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_34508_1577# 0
C343 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00205f
C344 swmatrix_Tgate_6.gated_control BUS[6] 0.86843f
C345 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_4921_1539# 0.0097f
C346 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C347 a_52860_1580# a_53228_2122# 0.00294f
C348 a_53376_2122# a_53580_2122# 0.01151f
C349 a_50912_2122# a_50764_2122# 0
C350 a_52392_1562# a_51256_2002# 0
C351 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C352 a_57396_1577# BUS[10] 0
C353 a_9900_2122# enable 0.00368f
C354 swmatrix_Tgate_3.gated_control PHI_1 0.01086f
C355 a_57356_2122# BUS[10] 0
C356 a_7084_2122# enable 0.00101f
C357 ShiftReg_row_10_2$1_0.Q[8] PHI_2 0.63578f
C358 a_40748_1577# PHI_2 0
C359 a_6248_1562# PHI_2 0.02762f
C360 swmatrix_Tgate_8.gated_control swmatrix_Tgate_4.gated_control 0.01259f
C361 a_49928_1562# swmatrix_Tgate_1.gated_control 0.01486f
C362 a_15788_2122# BUS[3] 0
C363 a_13816_2002# BUS[3] 0.0117f
C364 a_40380_1580# PHI_1 0.01277f
C365 a_40748_1577# BUS[7] 0
C366 a_39912_1562# PHI_1 0.01733f
C367 PHI_2 BUS[8] 0.11252f
C368 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C369 a_47136_2122# swmatrix_Tgate_3.gated_control 0.01553f
C370 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C371 a_9696_2122# vdd 0.55944f
C372 a_44672_2122# swmatrix_Tgate_3.gated_control 0.01496f
C373 a_1336_2002# enable 0.05124f
C374 a_7232_2122# vdd 0.56482f
C375 a_38776_2002# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C376 a_59468_2122# PHI_1 0.00164f
C377 swmatrix_Tgate_2.gated_control a_59468_1577# 0
C378 a_57496_2002# PHI_1 0.01314f
C379 ShiftReg_row_10_2$1_0.Q[6] a_36121_1539# 0.00241f
C380 a_28620_2122# PHI_2 0.00422f
C381 swmatrix_Tgate_1.gated_control a_56636_1580# 0
C382 a_56168_1562# a_57496_2002# 0.02403f
C383 a_25804_2122# PHI_2 0
C384 a_61081_1539# PHI_2 0
C385 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C386 a_3660_2122# PHI_1 0.00477f
C387 a_52860_1580# a_53720_2002# 0.00888f
C388 a_53376_2122# a_53228_2122# 0
C389 a_52392_1562# a_53720_2002# 0.02403f
C390 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_7.gated_control 0.23535f
C391 a_56168_1562# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C392 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_48601_1539# 0.0097f
C393 a_52392_1562# a_50396_1580# 0
C394 a_21660_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C395 d_out pin 0.01249f
C396 a_50912_2122# a_51256_2002# 0.57845f
C397 a_21192_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C398 a_59820_2122# BUS[10] 0.00104f
C399 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C400 a_9548_2122# enable 0.00101f
C401 ShiftReg_row_10_2$1_0.Q[3] a_20056_2002# 0.00242f
C402 a_57004_2122# BUS[10] 0
C403 a_49928_1562# PHI_1 0.70141f
C404 a_7576_2002# enable 0.05124f
C405 a_44524_1577# PHI_2 0
C406 a_41140_1577# PHI_2 0
C407 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C408 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C409 a_16280_2002# BUS[3] 0.01161f
C410 swmatrix_Tgate_9.gated_control D_in 0.17646f
C411 a_12488_1562# swmatrix_Tgate_4.gated_control 0.01486f
C412 a_12956_1580# BUS[3] 0.00688f
C413 a_40896_2122# PHI_1 0.01804f
C414 swmatrix_Tgate_4.gated_control PHI_2 0.31095f
C415 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C416 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C417 a_38432_2122# PHI_1 0.01882f
C418 a_41140_1577# BUS[7] 0
C419 a_26296_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C420 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C421 ShiftReg_row_10_2$1_0.Q[1] ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C422 a_41240_2002# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C423 swmatrix_Tgate_2.gated_control a_59860_1577# 0
C424 a_37916_1580# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C425 a_59960_2002# PHI_1 0.01261f
C426 a_56636_1580# PHI_1 0.0533f
C427 a_13676_2122# vdd 0.01506f
C428 a_28268_2122# PHI_2 0
C429 a_56168_1562# a_56636_1580# 0.30528f
C430 a_26296_2002# PHI_2 0.03207f
C431 a_59468_1577# PHI_2 0
C432 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN D_in 0
C433 a_3308_2122# PHI_1 0.00164f
C434 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C435 a_53376_2122# a_53720_2002# 0.57845f
C436 a_52392_1562# a_52860_1580# 0.30528f
C437 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_11161_1539# 0.0097f
C438 a_22176_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C439 ShiftReg_row_10_2$1_0.Q[6] vdd 0.57779f
C440 a_50912_2122# a_50396_1580# 0.30053f
C441 a_10040_2002# enable 0.0522f
C442 a_59468_2122# BUS[10] 0
C443 swmatrix_Tgate_7.gated_control BUS[3] 0.00566f
C444 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[8] 0.01102f
C445 a_44916_1577# PHI_2 0
C446 a_6716_1580# enable 0.05108f
C447 a_57496_2002# BUS[10] 0.0117f
C448 ShiftReg_row_10_2$1_0.Q[3] a_19196_1580# 0.36203f
C449 a_44876_2122# PHI_2 0.00411f
C450 a_15420_1580# BUS[3] 0.01336f
C451 a_14952_1562# BUS[3] 0.02637f
C452 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[10] 1.21861f
C453 a_18728_1562# PHI_2 0.02762f
C454 a_11161_1539# enable 0.00398f
C455 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[8] 0.10774f
C456 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C457 swmatrix_Tgate_3.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C458 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_28760_2002# 0.00242f
C459 a_25436_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C460 swmatrix_Tgate_7.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C461 ShiftReg_row_10_2$1_0.Q[1] a_4921_1539# 0.00241f
C462 pin BUS[3] 11.0719f
C463 a_59100_1580# PHI_1 0.01277f
C464 a_40380_1580# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C465 a_58632_1562# PHI_1 0.01733f
C466 a_39912_1562# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C467 a_16140_2122# vdd 0.01506f
C468 a_13324_2122# vdd 0.00491f
C469 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_8.gated_control 0.23535f
C470 ShiftReg_row_10_2$1_0.Q[6] a_38284_1577# 0
C471 a_9180_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C472 a_28760_2002# PHI_2 0.03174f
C473 a_56168_1562# a_58632_1562# 0
C474 a_8712_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C475 a_25436_1580# PHI_2 0.03321f
C476 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C477 a_3800_2002# PHI_1 0.01261f
C478 a_3800_2002# a_3700_1577# 0
C479 a_2940_1580# a_3308_1577# 0.00194f
C480 a_59860_1577# PHI_2 0
C481 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_7.gated_control 0.22418f
C482 swmatrix_Tgate_9.gated_control swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88175f
C483 a_53376_2122# a_52860_1580# 0.30053f
C484 a_52392_1562# a_53376_2122# 0.07055f
C485 a_50912_2122# a_52392_1562# 0.00268f
C486 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C487 PHI_1 BUS[6] 0.09486f
C488 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C489 a_59960_2002# BUS[10] 0.01161f
C490 swmatrix_Tgate_2.gated_control BUS[9] 0.00566f
C491 a_56636_1580# BUS[10] 0.00688f
C492 a_47340_2122# PHI_2 0.00422f
C493 a_9180_1580# enable 0.05124f
C494 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C495 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_6.gated_control 0.33472f
C496 a_8712_1562# enable 0.08694f
C497 a_44524_2122# PHI_2 0
C498 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C499 a_15420_1580# a_15788_1577# 0.00194f
C500 a_16280_2002# a_16180_1577# 0
C501 a_6248_1562# swmatrix_Tgate_9.gated_control 0.00493f
C502 a_15936_2122# BUS[3] 0.01571f
C503 ShiftReg_row_10_2$1_0.Q[3] enable 0.513f
C504 a_13472_2122# BUS[3] 0.0191f
C505 a_9548_1577# enable 0.0022f
C506 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C507 ShiftReg_row_10_2$1_0.Q[4] pin 0.01491f
C508 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_27900_1580# 0.36162f
C509 a_27432_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C510 a_476_1580# a_844_1577# 0.00194f
C511 a_59616_2122# PHI_1 0.01804f
C512 a_40896_2122# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C513 swmatrix_Tgate_6.gated_control PHI_2 0.31095f
C514 a_38432_2122# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C515 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C516 a_15788_2122# vdd 0.00491f
C517 a_57152_2122# PHI_1 0.01882f
C518 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C519 a_13816_2002# vdd 0.32603f
C520 a_8_1562# pin 0
C521 a_9696_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C522 a_27900_1580# PHI_2 0.07395f
C523 a_56168_1562# a_57152_2122# 0.07055f
C524 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C525 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C526 a_3456_2122# a_3308_1577# 0
C527 a_2940_1580# PHI_1 0.01277f
C528 a_27432_1562# PHI_2 0.60119f
C529 a_19564_1577# swmatrix_Tgate_7.gated_control 0
C530 ShiftReg_row_10_2$1_0.Q[4] a_24968_1562# 0.16779f
C531 a_13324_1577# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C532 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C533 a_32396_2122# vdd 0.01506f
C534 a_59100_1580# BUS[10] 0.01336f
C535 a_9696_2122# enable 0.11443f
C536 a_7232_2122# enable 0.11055f
C537 a_15936_2122# a_15788_1577# 0
C538 a_58632_1562# BUS[10] 0.02637f
C539 a_46988_2122# PHI_2 0
C540 ShiftReg_row_10_2$1_0.Q[3] a_19712_2122# 0.01552f
C541 a_7084_1577# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C542 a_45016_2002# PHI_2 0.03207f
C543 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_37448_1562# 0
C544 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C545 a_13324_1577# enable 0.0022f
C546 ShiftReg_row_10_2$1_0.Q[8] BUS[8] 0.01695f
C547 PHI_2 BUS[9] 0.11252f
C548 swmatrix_Tgate_5.gated_control a_29881_1539# 0.00113f
C549 a_31208_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C550 ShiftReg_row_10_2$1_0.Q[9] vdd 0.57779f
C551 a_9940_1577# enable 0.00579f
C552 a_28760_2002# ShiftReg_row_10_2$1_0.Q[5] 0.25874f
C553 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_28416_2122# 0.01536f
C554 ShiftReg_row_10_2$1_0.Q[9] ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C555 a_16180_1577# pin 0
C556 ShiftReg_row_10_2$1_0.Q[1] a_7084_1577# 0
C557 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_53228_1577# 0
C558 a_25952_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C559 ShiftReg_row_10_2$1_0.Q[1] PHI_1 0.05798f
C560 a_37448_1562# PHI_2 0.02762f
C561 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[9] 1.21861f
C562 a_16280_2002# vdd 0.32887f
C563 a_29881_1539# enable 0.00398f
C564 a_12956_1580# vdd 0.42253f
C565 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_8.gated_control 0.22418f
C566 swmatrix_Tgate_1.gated_control swmatrix_Tgate_2.gated_control 0.01259f
C567 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C568 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C569 a_28416_2122# PHI_2 0.04011f
C570 a_37448_1562# BUS[7] 0.0057f
C571 a_3456_2122# a_3700_1577# 0.01595f
C572 a_4921_1539# PHI_2 0
C573 a_3456_2122# PHI_1 0.01804f
C574 a_25952_2122# PHI_2 0.04895f
C575 a_19956_1577# swmatrix_Tgate_7.gated_control 0
C576 a_19916_2122# swmatrix_Tgate_7.gated_control 0
C577 a_34860_2122# vdd 0.01506f
C578 a_13716_1577# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C579 a_32044_2122# vdd 0.00491f
C580 a_8_1562# BUS[1] 0.00686f
C581 a_59616_2122# BUS[10] 0.01571f
C582 a_7476_1577# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C583 a_47480_2002# PHI_2 0.03174f
C584 a_57152_2122# BUS[10] 0.0191f
C585 a_15936_2122# a_16180_1577# 0.01595f
C586 a_44156_1580# PHI_2 0.03321f
C587 a_44524_1577# BUS[8] 0
C588 a_13716_1577# enable 0.00577f
C589 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_6.gated_control 0.17277f
C590 swmatrix_Tgate_5.gated_control a_28268_1577# 0
C591 a_13676_2122# enable 0.00368f
C592 a_27900_1580# ShiftReg_row_10_2$1_0.Q[5] 0.00101f
C593 a_19956_1577# pin 0
C594 a_25436_1580# a_25804_1577# 0.00194f
C595 a_27432_1562# ShiftReg_row_10_2$1_0.Q[5] 0.00225f
C596 a_26296_2002# a_26196_1577# 0
C597 ShiftReg_row_10_2$1_0.Q[9] a_54841_1539# 0.00241f
C598 a_26296_2002# a_26156_2122# 0.00109f
C599 swmatrix_Tgate_7.gated_control vdd 1.84761f
C600 a_29881_1539# BUS[5] 0
C601 ShiftReg_row_10_2$1_0.Q[6] enable 0.513f
C602 swmatrix_Tgate_2.gated_control PHI_1 0.00908f
C603 a_40380_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C604 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_0.gated_control 0.23535f
C605 a_28268_1577# enable 0.0022f
C606 a_7084_1577# swmatrix_Tgate_8.gated_control 0
C607 a_15420_1580# vdd 0.42496f
C608 ShiftReg_row_10_2$1_0.Q[2] a_12488_1562# 0.16779f
C609 a_56168_1562# swmatrix_Tgate_2.gated_control 0.01486f
C610 a_39912_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C611 a_14952_1562# vdd 1.0427f
C612 ShiftReg_row_10_2$1_0.Q[7] pin 0.01491f
C613 ShiftReg_row_10_2$1_0.Q[6] a_38776_2002# 0.00242f
C614 ShiftReg_row_10_2$1_0.Q[2] PHI_2 0.63578f
C615 swmatrix_Tgate_8.gated_control PHI_1 0.01086f
C616 a_3308_1577# PHI_2 0
C617 a_22380_2122# swmatrix_Tgate_7.gated_control 0
C618 swmatrix_Tgate_1.gated_control PHI_2 0.31095f
C619 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C620 a_34508_2122# vdd 0.00491f
C621 a_476_1580# pin 0.00137f
C622 swmatrix_Tgate_7.gated_control BUS[4] 0.86843f
C623 a_32536_2002# vdd 0.32603f
C624 vdd pin 10.3425f
C625 a_46620_1580# PHI_2 0.07395f
C626 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[9] 0
C627 a_45016_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C628 a_46152_1562# PHI_2 0.60119f
C629 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C630 swmatrix_Tgate_5.gated_control a_32044_1577# 0
C631 swmatrix_Tgate_5.gated_control a_28660_1577# 0
C632 a_44916_1577# BUS[8] 0
C633 swmatrix_Tgate_1.gated_control swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C634 a_16140_2122# enable 0.00368f
C635 a_13324_2122# enable 0.00101f
C636 a_44876_2122# BUS[8] 0
C637 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C638 a_51116_2122# vdd 0.01506f
C639 a_28416_2122# ShiftReg_row_10_2$1_0.Q[5] 0.11433f
C640 a_24968_1562# vdd 1.00067f
C641 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C642 a_28268_1577# BUS[5] 0
C643 pin BUS[4] 11.0719f
C644 a_40896_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C645 a_32044_1577# enable 0.0022f
C646 a_28660_1577# enable 0.00579f
C647 a_15936_2122# vdd 0.55944f
C648 a_7476_1577# swmatrix_Tgate_8.gated_control 0
C649 a_13472_2122# vdd 0.56482f
C650 a_7084_1577# PHI_2 0
C651 a_7436_2122# swmatrix_Tgate_8.gated_control 0
C652 a_3700_1577# PHI_2 0
C653 ShiftReg_row_10_2$1_0.Q[6] a_37916_1580# 0.36203f
C654 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C655 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C656 a_12488_1562# PHI_1 0.70141f
C657 PHI_1 PHI_2 24.2698f
C658 a_34900_1577# pin 0
C659 a_992_2122# PHI_2 0.04895f
C660 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C661 a_48601_1539# enable 0.00398f
C662 a_56168_1562# PHI_2 0.02762f
C663 a_35000_2002# vdd 0.32887f
C664 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[8] 1.21861f
C665 a_20056_2002# swmatrix_Tgate_7.gated_control 0.01121f
C666 PHI_1 BUS[7] 0.09486f
C667 a_31676_1580# vdd 0.42253f
C668 swmatrix_Tgate_2.gated_control BUS[10] 0.86843f
C669 a_2472_1562# pin 0.00127f
C670 a_13816_2002# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C671 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_47480_2002# 0.00242f
C672 a_47136_2122# PHI_2 0.04011f
C673 a_44156_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C674 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C675 a_844_1577# enable 0.0022f
C676 a_44672_2122# PHI_2 0.04895f
C677 a_7576_2002# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C678 a_15788_2122# enable 0.00101f
C679 a_53580_2122# vdd 0.01506f
C680 a_47340_2122# BUS[8] 0.00104f
C681 a_50764_2122# vdd 0.00491f
C682 vdd BUS[1] 0.56719f
C683 a_13816_2002# enable 0.05124f
C684 a_44524_2122# BUS[8] 0
C685 ShiftReg_row_10_2$1_0.Q[9] a_57004_1577# 0
C686 a_476_1580# BUS[1] 0.00598f
C687 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C688 a_28760_2002# a_28620_2122# 0.00109f
C689 a_18728_1562# swmatrix_Tgate_4.gated_control 0.00493f
C690 a_31208_1562# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C691 a_20056_2002# pin 0.00146f
C692 a_25952_2122# a_25804_1577# 0
C693 a_25436_1580# a_25804_2122# 0.00294f
C694 ShiftReg_row_10_2$1_0.Q[1] a_7576_2002# 0.00242f
C695 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_0.gated_control 0.22418f
C696 a_28660_1577# BUS[5] 0
C697 a_32436_1577# enable 0.00577f
C698 a_32396_2122# enable 0.00368f
C699 a_9900_2122# swmatrix_Tgate_8.gated_control 0
C700 a_7476_1577# PHI_2 0
C701 a_44524_1577# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C702 a_34140_1580# a_34508_1577# 0.00194f
C703 a_7436_2122# PHI_2 0.00411f
C704 a_38676_1577# pin 0
C705 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_1.gated_control 0.33472f
C706 a_35000_2002# a_34900_1577# 0
C707 swmatrix_Tgate_9.gated_control a_4921_1539# 0.00113f
C708 swmatrix_Tgate_0.gated_control vdd 1.84761f
C709 a_6248_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C710 a_22520_2002# swmatrix_Tgate_7.gated_control 0.01014f
C711 ShiftReg_row_10_2$1_0.Q[9] enable 0.513f
C712 a_46988_1577# enable 0.0022f
C713 a_19196_1580# swmatrix_Tgate_7.gated_control 0.00804f
C714 a_34140_1580# vdd 0.42496f
C715 a_33672_1562# vdd 1.0427f
C716 a_16280_2002# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C717 a_12956_1580# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C718 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C719 a_10040_2002# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C720 a_844_2122# PHI_2 0
C721 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_46620_1580# 0.36162f
C722 a_46152_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C723 a_6716_1580# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C724 a_1236_1577# enable 0.00577f
C725 a_46988_2122# BUS[8] 0
C726 a_16280_2002# enable 0.0522f
C727 a_53228_2122# vdd 0.00491f
C728 PHI_2 BUS[10] 0.11252f
C729 a_12956_1580# enable 0.05108f
C730 a_45016_2002# BUS[8] 0.0117f
C731 a_51256_2002# vdd 0.32603f
C732 a_2472_1562# BUS[1] 0.02735f
C733 ShiftReg_row_10_2$1_0.Q[5] PHI_1 0.05798f
C734 a_25952_2122# a_26196_1577# 0.01595f
C735 a_22520_2002# pin 0
C736 a_19196_1580# pin 0
C737 a_25952_2122# a_26156_2122# 0.01151f
C738 a_25436_1580# a_26296_2002# 0.00888f
C739 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[6] 0.10774f
C740 ShiftReg_row_10_2$1_0.Q[1] a_6716_1580# 0.36203f
C741 a_38284_1577# swmatrix_Tgate_0.gated_control 0
C742 ShiftReg_row_10_2$1_0.Q[7] a_43688_1562# 0.16779f
C743 a_34860_2122# enable 0.00368f
C744 a_32044_2122# enable 0.00101f
C745 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[1] 0.10851f
C746 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C747 a_9900_2122# PHI_2 0.00422f
C748 a_34656_2122# a_34508_1577# 0
C749 ShiftReg_row_10_2$1_0.Q[6] a_38432_2122# 0.01552f
C750 a_7576_2002# swmatrix_Tgate_8.gated_control 0.01121f
C751 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_56168_1562# 0
C752 swmatrix_Tgate_7.gated_control swmatrix_Tgate_5.gated_control 0.01259f
C753 a_44916_1577# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C754 a_7084_2122# PHI_2 0
C755 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C756 a_992_2122# D_in 0.01538f
C757 PHI_1 D_in 0.0221f
C758 a_43688_1562# vdd 1.00067f
C759 swmatrix_Tgate_7.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C760 swmatrix_Tgate_9.gated_control a_3308_1577# 0
C761 a_50764_1577# enable 0.0022f
C762 a_21660_1580# swmatrix_Tgate_7.gated_control 0.00668f
C763 a_49928_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C764 swmatrix_Tgate_3.gated_control a_48601_1539# 0.00113f
C765 a_47380_1577# enable 0.00579f
C766 a_34656_2122# vdd 0.55944f
C767 a_21192_1562# swmatrix_Tgate_7.gated_control 0.00985f
C768 a_47480_2002# ShiftReg_row_10_2$1_0.Q[8] 0.25874f
C769 a_15420_1580# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C770 a_32192_2122# vdd 0.56482f
C771 a_14952_1562# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C772 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_47136_2122# 0.01536f
C773 swmatrix_Tgate_7.gated_control enable 0.50846f
C774 ShiftReg_row_10_2$1_0.Q[3] ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C775 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C776 a_53620_1577# pin 0
C777 a_9180_1580# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C778 a_1336_2002# PHI_2 0.03207f
C779 a_44672_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C780 a_8712_1562# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C781 swmatrix_Tgate_5.gated_control pin 1.23291f
C782 a_47480_2002# BUS[8] 0.01161f
C783 a_15420_1580# enable 0.05124f
C784 a_14952_1562# enable 0.08694f
C785 a_53720_2002# vdd 0.32887f
C786 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[7] 1.21861f
C787 a_44156_1580# BUS[8] 0.00688f
C788 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C789 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C790 a_50396_1580# vdd 0.42253f
C791 a_28416_2122# a_28620_2122# 0.01151f
C792 a_27900_1580# a_28268_2122# 0.00294f
C793 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C794 a_21660_1580# pin 0.00113f
C795 a_25952_2122# a_25804_2122# 0
C796 a_21192_1562# pin 0.00138f
C797 a_27432_1562# a_26296_2002# 0
C798 a_38676_1577# swmatrix_Tgate_0.gated_control 0
C799 a_34508_2122# enable 0.00101f
C800 a_32536_2002# enable 0.05124f
C801 enable pin 1.18246f
C802 a_38636_2122# swmatrix_Tgate_0.gated_control 0
C803 a_10040_2002# swmatrix_Tgate_8.gated_control 0.01014f
C804 a_1196_2122# BUS[1] 0.00102f
C805 a_6716_1580# swmatrix_Tgate_8.gated_control 0.00804f
C806 a_9548_2122# PHI_2 0
C807 a_7576_2002# PHI_2 0.03207f
C808 swmatrix_Tgate_9.gated_control a_7084_1577# 0
C809 a_34656_2122# a_34900_1577# 0.01595f
C810 a_24968_1562# swmatrix_Tgate_5.gated_control 0.01486f
C811 a_38776_2002# pin 0.00146f
C812 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C813 swmatrix_Tgate_9.gated_control a_3700_1577# 0
C814 a_992_2122# swmatrix_Tgate_9.gated_control 0.01391f
C815 swmatrix_Tgate_9.gated_control PHI_1 0.01082f
C816 a_51156_1577# enable 0.00577f
C817 a_22176_2122# swmatrix_Tgate_7.gated_control 0.01553f
C818 ShiftReg_row_10_2$1_0.Q[8] swmatrix_Tgate_1.gated_control 0.17277f
C819 a_51116_2122# enable 0.00368f
C820 swmatrix_Tgate_8.gated_control a_11161_1539# 0.00113f
C821 a_19712_2122# swmatrix_Tgate_7.gated_control 0.01496f
C822 swmatrix_Tgate_3.gated_control a_46988_1577# 0
C823 a_12488_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C824 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C825 a_15936_2122# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C826 a_13472_2122# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C827 a_46620_1580# ShiftReg_row_10_2$1_0.Q[8] 0.00101f
C828 a_24968_1562# enable 0.08752f
C829 a_44156_1580# a_44524_1577# 0.00194f
C830 a_57396_1577# pin 0
C831 swmatrix_Tgate_1.gated_control BUS[8] 0.00566f
C832 a_45016_2002# a_44916_1577# 0
C833 a_46152_1562# ShiftReg_row_10_2$1_0.Q[8] 0.00225f
C834 a_45016_2002# a_44876_2122# 0.00109f
C835 a_9696_2122# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C836 a_7232_2122# swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C837 a_46620_1580# BUS[8] 0.01336f
C838 a_15936_2122# enable 0.11443f
C839 a_31208_1562# a_32536_2002# 0.02403f
C840 a_31208_1562# pin 0
C841 swmatrix_Tgate_5.gated_control a_31676_1580# 0
C842 a_13472_2122# enable 0.11055f
C843 a_52860_1580# vdd 0.42496f
C844 a_46152_1562# BUS[8] 0.02637f
C845 a_52392_1562# vdd 1.0427f
C846 a_28416_2122# a_28268_2122# 0
C847 a_27900_1580# a_28760_2002# 0.00888f
C848 ShiftReg_row_10_2$1_0.Q[9] a_57496_2002# 0.00242f
C849 a_22176_2122# pin 0.00251f
C850 ShiftReg_row_10_2$1_0.Q[6] BUS[6] 0.01695f
C851 a_27432_1562# a_28760_2002# 0.02403f
C852 a_19712_2122# pin 0.00138f
C853 a_992_2122# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C854 a_26156_2122# PHI_1 0.00534f
C855 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_23641_1539# 0.0097f
C856 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0.0011f
C857 a_25952_2122# a_26296_2002# 0.57845f
C858 a_27432_1562# a_25436_1580# 0
C859 pin BUS[5] 11.0719f
C860 ShiftReg_row_10_2$1_0.Q[1] a_7232_2122# 0.01552f
C861 a_41100_2122# swmatrix_Tgate_0.gated_control 0
C862 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C863 a_35000_2002# enable 0.0522f
C864 a_31676_1580# enable 0.05108f
C865 a_9180_1580# swmatrix_Tgate_8.gated_control 0.00668f
C866 a_8712_1562# swmatrix_Tgate_8.gated_control 0.00985f
C867 a_10040_2002# PHI_2 0.03174f
C868 a_41240_2002# pin 0
C869 a_45016_2002# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C870 a_6716_1580# PHI_2 0.03321f
C871 ShiftReg_row_10_2$1_0.Q[8] PHI_1 0.05798f
C872 a_37916_1580# pin 0
C873 swmatrix_Tgate_3.gated_control a_50764_1577# 0
C874 ShiftReg_row_10_2$1_0.Q[2] swmatrix_Tgate_4.gated_control 0.17277f
C875 a_6248_1562# PHI_1 0.70141f
C876 enable BUS[1] 0.21583f
C877 a_53580_2122# enable 0.00368f
C878 swmatrix_Tgate_3.gated_control a_47380_1577# 0
C879 swmatrix_Tgate_8.gated_control a_9548_1577# 0
C880 a_50764_2122# enable 0.00101f
C881 a_11161_1539# PHI_2 0
C882 PHI_1 BUS[8] 0.09486f
C883 a_24968_1562# BUS[5] 0.0057f
C884 a_47136_2122# ShiftReg_row_10_2$1_0.Q[8] 0.11433f
C885 a_1336_2002# D_in 0.00242f
C886 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C887 a_47136_2122# BUS[8] 0.01571f
C888 vdd BUS[2] 0.56053f
C889 a_53376_2122# vdd 0.55944f
C890 a_31208_1562# a_31676_1580# 0.30528f
C891 a_44672_2122# BUS[8] 0.0191f
C892 a_50912_2122# vdd 0.56482f
C893 swmatrix_Tgate_0.gated_control enable 0.50846f
C894 a_28416_2122# a_28760_2002# 0.57845f
C895 a_28620_2122# PHI_1 0.00477f
C896 ShiftReg_row_10_2$1_0.Q[9] a_56636_1580# 0.36203f
C897 a_25804_2122# PHI_1 0.00201f
C898 a_32044_1577# BUS[6] 0
C899 a_27432_1562# a_27900_1580# 0.30528f
C900 a_25952_2122# a_25436_1580# 0.30053f
C901 a_38776_2002# swmatrix_Tgate_0.gated_control 0.01121f
C902 swmatrix_Tgate_3.gated_control pin 1.23291f
C903 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[4] 0.01102f
C904 a_34140_1580# enable 0.05124f
C905 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[6] 1.21861f
C906 a_33672_1562# enable 0.08694f
C907 a_9696_2122# swmatrix_Tgate_8.gated_control 0.01553f
C908 a_9180_1580# PHI_2 0.07395f
C909 a_47480_2002# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C910 a_7232_2122# swmatrix_Tgate_8.gated_control 0.01496f
C911 a_17401_1539# BUS[3] 0
C912 a_40380_1580# pin 0.00113f
C913 a_44156_1580# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C914 a_39912_1562# pin 0.00138f
C915 a_8712_1562# PHI_2 0.60119f
C916 swmatrix_Tgate_8.gated_control a_13324_1577# 0
C917 ShiftReg_row_10_2$1_0.Q[3] PHI_2 0.63578f
C918 swmatrix_Tgate_8.gated_control a_9940_1577# 0
C919 a_53228_2122# enable 0.00101f
C920 a_9548_1577# PHI_2 0
C921 swmatrix_Tgate_4.gated_control PHI_1 0.01086f
C922 a_51256_2002# enable 0.05124f
C923 a_37448_1562# swmatrix_Tgate_6.gated_control 0.00493f
C924 a_47480_2002# a_47340_2122# 0.00109f
C925 a_44672_2122# a_44524_1577# 0
C926 a_57496_2002# pin 0.00146f
C927 a_44156_1580# a_44524_2122# 0.00294f
C928 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C929 a_1336_2002# swmatrix_Tgate_9.gated_control 0.01107f
C930 a_31208_1562# a_33672_1562# 0
C931 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C932 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C933 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[7] 0
C934 a_28416_2122# a_27900_1580# 0.30053f
C935 a_28268_2122# PHI_1 0.00164f
C936 a_52860_1580# a_53228_1577# 0.00194f
C937 a_43688_1562# enable 0.08752f
C938 a_27432_1562# a_28416_2122# 0.07055f
C939 a_53720_2002# a_53620_1577# 0
C940 a_26296_2002# PHI_1 0.01314f
C941 a_25952_2122# a_27432_1562# 0.00268f
C942 a_32436_1577# BUS[6] 0
C943 a_32396_2122# BUS[6] 0
C944 a_34656_2122# enable 0.11443f
C945 swmatrix_Tgate_1.gated_control swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C946 a_41240_2002# swmatrix_Tgate_0.gated_control 0.01014f
C947 a_37916_1580# swmatrix_Tgate_0.gated_control 0.00804f
C948 a_49928_1562# pin 0
C949 a_32192_2122# enable 0.11055f
C950 swmatrix_Tgate_5.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C951 a_40896_2122# pin 0.00251f
C952 a_9696_2122# PHI_2 0.04011f
C953 a_46620_1580# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C954 a_15788_1577# BUS[3] 0
C955 a_46152_1562# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C956 a_7232_2122# PHI_2 0.04895f
C957 a_44876_2122# PHI_1 0.00534f
C958 a_38432_2122# pin 0.00138f
C959 a_1336_2002# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C960 a_53720_2002# enable 0.0522f
C961 a_18728_1562# PHI_1 0.70141f
C962 a_13324_1577# PHI_2 0
C963 a_50396_1580# enable 0.05108f
C964 a_9940_1577# PHI_2 0
C965 a_61081_1539# BUS[10] 0
C966 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C967 a_44672_2122# a_44916_1577# 0.01595f
C968 a_59960_2002# pin 0
C969 a_44156_1580# a_45016_2002# 0.00888f
C970 a_56636_1580# pin 0
C971 a_44672_2122# a_44876_2122# 0.01151f
C972 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C973 a_29881_1539# PHI_2 0
C974 a_31208_1562# a_32192_2122# 0.07055f
C975 a_53376_2122# a_53228_1577# 0
C976 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[2] 0.01102f
C977 ShiftReg_row_10_2$1_0.Q[9] a_57152_2122# 0.01552f
C978 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C979 swmatrix_Tgate_0.gated_control swmatrix_Tgate_3.gated_control 0.01259f
C980 a_28760_2002# PHI_1 0.01261f
C981 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C982 a_34860_2122# BUS[6] 0.00104f
C983 a_25436_1580# PHI_1 0.0533f
C984 a_32044_2122# BUS[6] 0
C985 a_40380_1580# swmatrix_Tgate_0.gated_control 0.00668f
C986 a_3660_2122# BUS[1] 0.00101f
C987 a_39912_1562# swmatrix_Tgate_0.gated_control 0.00985f
C988 vdd d_out 0.40535f
C989 ShiftReg_row_10_2$1_0.Q[6] ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C990 a_47340_2122# PHI_1 0.00477f
C991 a_16180_1577# BUS[3] 0
C992 a_47136_2122# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C993 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q d_out 0.01102f
C994 a_6248_1562# a_7576_2002# 0.02403f
C995 a_44524_2122# PHI_1 0.00201f
C996 swmatrix_Tgate_9.gated_control a_6716_1580# 0
C997 a_44672_2122# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C998 a_52860_1580# enable 0.05124f
C999 a_52392_1562# enable 0.08694f
C1000 ShiftReg_row_10_2$1_0.Q[5] ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C1001 a_59468_1577# BUS[10] 0
C1002 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[5] 1.21861f
C1003 a_13716_1577# PHI_2 0
C1004 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_28268_1577# 0
C1005 a_13676_2122# PHI_2 0.00411f
C1006 a_46620_1580# a_46988_2122# 0.00294f
C1007 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1008 a_47136_2122# a_47340_2122# 0.01151f
C1009 swmatrix_Tgate_1.gated_control BUS[9] 0.86843f
C1010 a_59100_1580# pin 0.00113f
C1011 a_44672_2122# a_44524_2122# 0
C1012 a_46152_1562# a_45016_2002# 0
C1013 a_58632_1562# pin 0.00138f
C1014 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C1015 a_19564_1577# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1016 ShiftReg_row_10_2$1_0.Q[6] PHI_2 0.63578f
C1017 swmatrix_Tgate_6.gated_control PHI_1 0.01086f
C1018 a_28268_1577# PHI_2 0
C1019 a_3800_2002# pin 0
C1020 a_43688_1562# swmatrix_Tgate_3.gated_control 0.01486f
C1021 a_53376_2122# a_53620_1577# 0.01595f
C1022 a_34508_2122# BUS[6] 0
C1023 a_27900_1580# PHI_1 0.01277f
C1024 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C1025 pin BUS[6] 11.0719f
C1026 a_27432_1562# PHI_1 0.01733f
C1027 a_32536_2002# BUS[6] 0.0117f
C1028 a_40896_2122# swmatrix_Tgate_0.gated_control 0.01553f
C1029 a_38432_2122# swmatrix_Tgate_0.gated_control 0.01496f
C1030 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[2] 0
C1031 a_3308_2122# BUS[1] 0
C1032 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C1033 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[4] 0.10774f
C1034 a_46988_2122# PHI_1 0.00164f
C1035 a_45016_2002# PHI_1 0.01314f
C1036 a_6248_1562# a_6716_1580# 0.30528f
C1037 ShiftReg_row_10_2$1_0.Q[5] a_29881_1539# 0.00241f
C1038 swmatrix_Tgate_3.gated_control a_50396_1580# 0
C1039 a_16140_2122# PHI_2 0.00422f
C1040 enable BUS[2] 0.2115f
C1041 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1042 a_49928_1562# a_51256_2002# 0.02403f
C1043 a_53376_2122# enable 0.11443f
C1044 a_59860_1577# BUS[10] 0
C1045 a_50912_2122# enable 0.11055f
C1046 PHI_1 BUS[9] 0.09486f
C1047 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C1048 a_13324_2122# PHI_2 0
C1049 a_46620_1580# a_47480_2002# 0.00888f
C1050 a_47136_2122# a_46988_2122# 0
C1051 a_59616_2122# pin 0.00251f
C1052 a_46152_1562# a_47480_2002# 0.02403f
C1053 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_4.gated_control 0.23535f
C1054 a_15420_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1055 a_46152_1562# a_44156_1580# 0
C1056 a_57152_2122# pin 0.00138f
C1057 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_42361_1539# 0.0097f
C1058 a_14952_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1059 a_44672_2122# a_45016_2002# 0.57845f
C1060 a_19956_1577# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1061 a_32044_1577# PHI_2 0
C1062 vdd BUS[3] 0.56053f
C1063 a_37448_1562# PHI_1 0.70141f
C1064 a_28660_1577# PHI_2 0
C1065 a_2940_1580# pin 0.00108f
C1066 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_2.gated_control 0.17277f
C1067 a_28416_2122# PHI_1 0.01804f
C1068 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C1069 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C1070 a_35000_2002# BUS[6] 0.01161f
C1071 a_25952_2122# PHI_1 0.01882f
C1072 a_31676_1580# BUS[6] 0.00688f
C1073 a_48601_1539# PHI_2 0
C1074 a_3800_2002# BUS[1] 0.01037f
C1075 a_20056_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1076 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57452f
C1077 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN d_out 0.08537f
C1078 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C1079 a_47480_2002# PHI_1 0.01261f
C1080 a_44156_1580# PHI_1 0.0533f
C1081 a_844_1577# PHI_2 0
C1082 a_6248_1562# a_8712_1562# 0
C1083 swmatrix_Tgate_8.gated_control a_12956_1580# 0
C1084 a_49928_1562# a_50396_1580# 0.30528f
C1085 a_12488_1562# a_13816_2002# 0.02403f
C1086 a_15788_2122# PHI_2 0
C1087 a_13816_2002# PHI_2 0.03207f
C1088 ShiftReg_row_10_2$1_0.Q[1] pin 0.01507f
C1089 a_47136_2122# a_47480_2002# 0.57845f
C1090 a_46152_1562# a_46620_1580# 0.30528f
C1091 a_15936_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1092 a_44672_2122# a_44156_1580# 0.30053f
C1093 ShiftReg_row_10_2$1_0.Q[4] vdd 0.57779f
C1094 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[7] 0.01102f
C1095 a_32436_1577# PHI_2 0
C1096 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[4] 1.21861f
C1097 a_3456_2122# pin 0
C1098 swmatrix_Tgate_0.gated_control BUS[6] 0.00566f
C1099 a_32396_2122# PHI_2 0.00411f
C1100 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1101 ShiftReg_row_10_2$1_0.Q[2] PHI_1 0.05798f
C1102 a_8_1562# vdd 0.99867f
C1103 a_34140_1580# BUS[6] 0.01336f
C1104 a_8_1562# a_476_1580# 0.30528f
C1105 a_33672_1562# BUS[6] 0.02637f
C1106 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C1107 ShiftReg_row_10_2$1_0.Q[9] PHI_2 0.63578f
C1108 swmatrix_Tgate_1.gated_control PHI_1 0.01086f
C1109 a_46988_1577# PHI_2 0
C1110 a_2940_1580# BUS[1] 0.01251f
C1111 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_22520_2002# 0.00242f
C1112 a_19196_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1113 ShiftReg_row_10_2$1_0.Q[4] BUS[4] 0.01695f
C1114 a_56168_1562# swmatrix_Tgate_1.gated_control 0.00493f
C1115 a_46620_1580# PHI_1 0.01277f
C1116 a_1236_1577# PHI_2 0
C1117 a_46152_1562# PHI_1 0.01733f
C1118 a_6248_1562# a_7232_2122# 0.07055f
C1119 ShiftReg_row_10_2$1_0.Q[5] a_32044_1577# 0
C1120 a_12488_1562# a_12956_1580# 0.30528f
C1121 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C1122 a_49928_1562# a_52392_1562# 0
C1123 a_16280_2002# PHI_2 0.03174f
C1124 a_12956_1580# PHI_2 0.03321f
C1125 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1126 swmatrix_Tgate_2.gated_control pin 1.23291f
C1127 a_47136_2122# a_46620_1580# 0.30053f
C1128 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_4.gated_control 0.22418f
C1129 a_46152_1562# a_47136_2122# 0.07055f
C1130 a_44672_2122# a_46152_1562# 0.00268f
C1131 a_20056_2002# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1132 enable d_out 0.38669f
C1133 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_5.gated_control 0.33472f
C1134 swmatrix_Tgate_8.gated_control pin 1.23275f
C1135 a_34860_2122# PHI_2 0.00422f
C1136 a_32044_2122# PHI_2 0
C1137 ShiftReg_row_10_2$1_0.Q[1] BUS[1] 0.00756f
C1138 a_7576_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1139 a_34656_2122# BUS[6] 0.01571f
C1140 a_8_1562# a_2472_1562# 0
C1141 a_992_2122# PHI_1 0.01882f
C1142 a_32192_2122# BUS[6] 0.0191f
C1143 a_56168_1562# PHI_1 0.70141f
C1144 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_21660_1580# 0.36162f
C1145 a_37448_1562# swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1146 a_50764_1577# PHI_2 0
C1147 a_21192_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1148 a_47380_1577# PHI_2 0
C1149 a_3456_2122# BUS[1] 0.01882f
C1150 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1151 a_19564_1577# BUS[4] 0
C1152 a_47136_2122# PHI_1 0.01804f
C1153 a_8_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C1154 swmatrix_Tgate_7.gated_control PHI_2 0.31095f
C1155 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C1156 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C1157 a_844_1577# D_in 0
C1158 a_44672_2122# PHI_1 0.01882f
C1159 a_12488_1562# a_14952_1562# 0
C1160 a_50764_1577# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1161 a_49928_1562# a_50912_2122# 0.07055f
C1162 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C1163 a_15420_1580# PHI_2 0.07395f
C1164 a_14952_1562# PHI_2 0.60119f
C1165 a_13324_1577# swmatrix_Tgate_4.gated_control 0
C1166 ShiftReg_row_10_2$1_0.Q[3] a_18728_1562# 0.16779f
C1167 a_19916_2122# vdd 0.01506f
C1168 a_22520_2002# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C1169 a_19196_1580# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1170 a_12488_1562# pin 0
C1171 PHI_2 pin 0.12723f
C1172 a_34508_2122# PHI_2 0
C1173 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_31208_1562# 0
C1174 a_32536_2002# PHI_2 0.03207f
C1175 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_10040_2002# 0.00242f
C1176 a_6716_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1177 ShiftReg_row_10_2$1_0.Q[9] ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1178 ShiftReg_row_10_2$1_0.Q[7] vdd 0.57779f
C1179 a_7436_2122# PHI_1 0.00534f
C1180 swmatrix_Tgate_7.gated_control a_23641_1539# 0.00113f
C1181 a_24968_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C1182 pin BUS[7] 11.0719f
C1183 swmatrix_Tgate_8.gated_control BUS[1] 0.00492f
C1184 a_22520_2002# ShiftReg_row_10_2$1_0.Q[4] 0.25874f
C1185 ShiftReg_row_10_2$1_0.Q[8] ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C1186 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[5] 0
C1187 a_51156_1577# PHI_2 0
C1188 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_46988_1577# 0
C1189 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_22176_2122# 0.01536f
C1190 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[3] 1.21861f
C1191 a_19712_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C1192 a_51116_2122# PHI_2 0.00411f
C1193 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C1194 a_19956_1577# BUS[4] 0
C1195 a_476_1580# vdd 0.42254f
C1196 a_19916_2122# BUS[4] 0
C1197 a_992_2122# a_844_2122# 0
C1198 a_844_2122# PHI_1 0.00201f
C1199 a_24968_1562# PHI_2 0.02762f
C1200 a_17401_1539# enable 0.00398f
C1201 a_844_1577# swmatrix_Tgate_9.gated_control 0
C1202 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C1203 enable BUS[3] 0.2115f
C1204 PHI_1 BUS[10] 0.09486f
C1205 a_12488_1562# a_13472_2122# 0.07055f
C1206 a_51156_1577# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1207 a_15936_2122# PHI_2 0.04011f
C1208 a_13472_2122# PHI_2 0.04895f
C1209 swmatrix_Tgate_5.gated_control swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C1210 a_56168_1562# BUS[10] 0.0057f
C1211 a_13716_1577# swmatrix_Tgate_4.gated_control 0
C1212 a_13676_2122# swmatrix_Tgate_4.gated_control 0
C1213 a_22380_2122# vdd 0.01506f
C1214 a_19564_2122# vdd 0.00491f
C1215 a_21660_1580# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C1216 vdd BUS[4] 0.56053f
C1217 a_21192_1562# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C1218 a_35000_2002# PHI_2 0.03174f
C1219 a_31676_1580# PHI_2 0.03321f
C1220 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C1221 a_9900_2122# PHI_1 0.00477f
C1222 ShiftReg_row_10_2$1_0.Q[4] swmatrix_Tgate_5.gated_control 0.17277f
C1223 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_9180_1580# 0.36162f
C1224 a_7084_2122# PHI_1 0.00201f
C1225 a_8712_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1226 swmatrix_Tgate_7.gated_control a_22028_1577# 0
C1227 a_844_1577# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1228 ShiftReg_row_10_2$1_0.Q[8] a_48601_1539# 0.00241f
C1229 a_21660_1580# ShiftReg_row_10_2$1_0.Q[4] 0.00101f
C1230 ShiftReg_row_10_2$1_0.Q[2] ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C1231 a_53580_2122# PHI_2 0.00422f
C1232 a_20056_2002# a_19956_1577# 0
C1233 a_21192_1562# ShiftReg_row_10_2$1_0.Q[4] 0.00225f
C1234 a_50764_2122# PHI_2 0
C1235 PHI_2 BUS[1] 0.10474f
C1236 a_19196_1580# a_19564_1577# 0.00194f
C1237 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_9548_1577# 0
C1238 a_20056_2002# a_19916_2122# 0.00109f
C1239 a_22380_2122# BUS[4] 0.00104f
C1240 a_19564_2122# BUS[4] 0
C1241 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_6.gated_control 0.23535f
C1242 a_34140_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1243 ShiftReg_row_10_2$1_0.Q[4] enable 0.513f
C1244 a_2472_1562# vdd 1.04366f
C1245 a_48601_1539# BUS[8] 0
C1246 a_2472_1562# a_476_1580# 0
C1247 a_15788_1577# enable 0.0022f
C1248 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C1249 a_992_2122# a_1336_2002# 0.57845f
C1250 a_1336_2002# PHI_1 0.01314f
C1251 a_33672_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1252 a_1236_1577# swmatrix_Tgate_9.gated_control 0
C1253 ShiftReg_row_10_2$1_0.Q[5] pin 0.01491f
C1254 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1255 ShiftReg_row_10_2$1_0.Q[5] a_32536_2002# 0.00242f
C1256 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN d_out 0.00347f
C1257 swmatrix_Tgate_0.gated_control PHI_2 0.31095f
C1258 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34499f
C1259 a_8_1562# enable 0.08666f
C1260 a_16140_2122# swmatrix_Tgate_4.gated_control 0
C1261 a_22028_2122# vdd 0.00491f
C1262 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C1263 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C1264 a_476_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1265 a_20056_2002# vdd 0.32603f
C1266 a_22176_2122# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C1267 a_19712_2122# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1268 a_34140_1580# PHI_2 0.07395f
C1269 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C1270 swmatrix_Tgate_0.gated_control BUS[7] 0.86843f
C1271 D_in pin 0.00593f
C1272 a_33672_1562# PHI_2 0.60119f
C1273 a_38776_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1274 a_10040_2002# ShiftReg_row_10_2$1_0.Q[2] 0.25874f
C1275 a_9548_2122# PHI_1 0.00164f
C1276 swmatrix_Tgate_7.gated_control a_25804_1577# 0
C1277 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_9696_2122# 0.01536f
C1278 a_7576_2002# PHI_1 0.01314f
C1279 a_7232_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C1280 swmatrix_Tgate_7.gated_control a_22420_1577# 0
C1281 a_1236_1577# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1282 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C1283 a_38636_2122# vdd 0.01506f
C1284 a_22176_2122# ShiftReg_row_10_2$1_0.Q[4] 0.11433f
C1285 ShiftReg_row_10_2$1_0.Q[2] a_11161_1539# 0.00241f
C1286 a_53228_2122# PHI_2 0
C1287 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C1288 a_51256_2002# PHI_2 0.03207f
C1289 a_22028_2122# BUS[4] 0
C1290 a_20056_2002# BUS[4] 0.0117f
C1291 a_59960_2002# d_out 0.25874f
C1292 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42601f
C1293 a_19564_1577# enable 0.0022f
C1294 a_34656_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1295 a_46988_1577# BUS[8] 0
C1296 a_16180_1577# enable 0.00579f
C1297 a_22420_1577# pin 0
C1298 ShiftReg_row_10_2$1_0.Q[5] a_31676_1580# 0.36203f
C1299 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[2] 1.21861f
C1300 a_51256_2002# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1301 a_1196_2122# vdd 0.01506f
C1302 a_43688_1562# PHI_2 0.02762f
C1303 a_2472_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1304 a_36121_1539# enable 0.00398f
C1305 a_22520_2002# vdd 0.32887f
C1306 a_13816_2002# swmatrix_Tgate_4.gated_control 0.01121f
C1307 a_19196_1580# vdd 0.42253f
C1308 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_41240_2002# 0.00242f
C1309 a_34656_2122# PHI_2 0.04011f
C1310 a_32192_2122# PHI_2 0.04895f
C1311 swmatrix_Tgate_9.gated_control pin 1.22292f
C1312 a_9180_1580# ShiftReg_row_10_2$1_0.Q[2] 0.00101f
C1313 a_37916_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1314 a_7576_2002# a_7476_1577# 0
C1315 a_8712_1562# ShiftReg_row_10_2$1_0.Q[2] 0.00225f
C1316 a_6716_1580# a_7084_1577# 0.00194f
C1317 a_7576_2002# a_7436_2122# 0.00109f
C1318 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C1319 a_10040_2002# PHI_1 0.01261f
C1320 a_41100_2122# vdd 0.01506f
C1321 a_6716_1580# PHI_1 0.0533f
C1322 a_38284_2122# vdd 0.00491f
C1323 a_22520_2002# a_22380_2122# 0.00109f
C1324 ShiftReg_row_10_2$1_0.Q[8] a_50764_1577# 0
C1325 a_19712_2122# a_19564_1577# 0
C1326 a_53720_2002# PHI_2 0.03174f
C1327 D_in BUS[1] 0.00379f
C1328 a_19196_1580# a_19564_2122# 0.00294f
C1329 a_50396_1580# PHI_2 0.03321f
C1330 a_22520_2002# BUS[4] 0.01161f
C1331 a_59100_1580# d_out 0.00101f
C1332 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_6.gated_control 0.22418f
C1333 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C1334 a_19956_1577# enable 0.00577f
C1335 a_19196_1580# BUS[4] 0.00688f
C1336 a_58632_1562# d_out 0.00225f
C1337 a_19916_2122# enable 0.00368f
C1338 a_47380_1577# BUS[8] 0
C1339 a_27900_1580# a_28268_1577# 0.00194f
C1340 a_53720_2002# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C1341 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_3.gated_control 0.33472f
C1342 a_28760_2002# a_28660_1577# 0
C1343 a_26196_1577# pin 0
C1344 swmatrix_Tgate_5.gated_control vdd 1.84761f
C1345 a_50396_1580# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1346 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57323f
C1347 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1348 ShiftReg_row_10_2$1_0.Q[7] enable 0.513f
C1349 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C1350 a_16280_2002# swmatrix_Tgate_4.gated_control 0.01014f
C1351 a_34508_1577# enable 0.0022f
C1352 a_21660_1580# vdd 0.42496f
C1353 a_12956_1580# swmatrix_Tgate_4.gated_control 0.00804f
C1354 a_21192_1562# vdd 1.0427f
C1355 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_40380_1580# 0.36162f
C1356 ShiftReg_row_10_2$1_0.Q[8] pin 0.01491f
C1357 a_39912_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1358 a_6248_1562# pin 0
C1359 vdd enable 4.10346f
C1360 a_9696_2122# ShiftReg_row_10_2$1_0.Q[2] 0.11433f
C1361 a_476_1580# enable 0.05107f
C1362 a_9180_1580# PHI_1 0.01277f
C1363 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C1364 a_40748_2122# vdd 0.00491f
C1365 pin BUS[8] 11.0719f
C1366 a_8712_1562# PHI_1 0.01733f
C1367 ShiftReg_row_10_2$1_0.Q[2] a_13324_1577# 0
C1368 swmatrix_Tgate_5.gated_control BUS[4] 0.00566f
C1369 swmatrix_Tgate_8.gated_control BUS[2] 0.86843f
C1370 a_38776_2002# vdd 0.32603f
C1371 a_52860_1580# PHI_2 0.07395f
C1372 a_52392_1562# PHI_2 0.60119f
C1373 a_19712_2122# a_19956_1577# 0.01595f
C1374 ShiftReg_row_10_2$1_0.Q[3] PHI_1 0.05798f
C1375 a_19712_2122# a_19916_2122# 0.01151f
C1376 a_19196_1580# a_20056_2002# 0.00888f
C1377 swmatrix_Tgate_9.gated_control BUS[1] 0.88604f
C1378 a_21660_1580# BUS[4] 0.01336f
C1379 a_22380_2122# enable 0.00368f
C1380 a_21192_1562# BUS[4] 0.02637f
C1381 a_32044_1577# swmatrix_Tgate_6.gated_control 0
C1382 a_59616_2122# d_out 0.11433f
C1383 ShiftReg_row_10_2$1_0.Q[6] a_37448_1562# 0.16779f
C1384 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[9] 0.10774f
C1385 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C1386 a_19564_2122# enable 0.00101f
C1387 a_57356_2122# vdd 0.01506f
C1388 swmatrix_Tgate_6.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C1389 enable BUS[4] 0.2115f
C1390 a_28416_2122# a_28268_1577# 0
C1391 ShiftReg_row_10_2$1_0.Q[5] a_32192_2122# 0.01552f
C1392 a_52860_1580# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C1393 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_49928_1562# 0
C1394 swmatrix_Tgate_4.gated_control swmatrix_Tgate_7.gated_control 0.01259f
C1395 a_52392_1562# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C1396 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C1397 a_31208_1562# vdd 1.00067f
C1398 a_38284_1577# enable 0.0022f
C1399 a_15420_1580# swmatrix_Tgate_4.gated_control 0.00668f
C1400 a_34900_1577# enable 0.00579f
C1401 a_43688_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C1402 swmatrix_Tgate_0.gated_control a_42361_1539# 0.00113f
C1403 a_14952_1562# swmatrix_Tgate_4.gated_control 0.00985f
C1404 a_22176_2122# vdd 0.55944f
C1405 a_41240_2002# ShiftReg_row_10_2$1_0.Q[7] 0.25874f
C1406 a_19712_2122# vdd 0.56482f
C1407 vdd BUS[5] 0.56053f
C1408 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_40896_2122# 0.01536f
C1409 a_41140_1577# pin 0
C1410 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN BUS[1] 1.21878f
C1411 a_38432_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C1412 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C1413 a_10040_2002# a_9900_2122# 0.00109f
C1414 a_2472_1562# enable 0.08694f
C1415 a_9696_2122# PHI_1 0.01804f
C1416 a_7232_2122# a_7084_1577# 0
C1417 a_6716_1580# a_7084_2122# 0.00294f
C1418 swmatrix_Tgate_4.gated_control pin 1.23291f
C1419 a_54841_1539# enable 0.00398f
C1420 a_7232_2122# PHI_1 0.01882f
C1421 a_41240_2002# vdd 0.32887f
C1422 a_37916_1580# vdd 0.42253f
C1423 PHI_2 BUS[2] 0.11252f
C1424 a_53376_2122# PHI_2 0.04011f
C1425 a_22176_2122# a_22380_2122# 0.01151f
C1426 a_21660_1580# a_22028_2122# 0.00294f
C1427 a_50912_2122# PHI_2 0.04895f
C1428 a_19712_2122# a_19564_2122# 0
C1429 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C1430 a_21192_1562# a_20056_2002# 0
C1431 a_22176_2122# BUS[4] 0.01571f
C1432 a_32436_1577# swmatrix_Tgate_6.gated_control 0
C1433 a_19712_2122# BUS[4] 0.0191f
C1434 a_32396_2122# swmatrix_Tgate_6.gated_control 0
C1435 a_22028_2122# enable 0.00101f
C1436 a_20056_2002# enable 0.05124f
C1437 a_59820_2122# vdd 0.01506f
C1438 a_57004_2122# vdd 0.00491f
C1439 a_18728_1562# swmatrix_Tgate_7.gated_control 0.01486f
C1440 a_28416_2122# a_28660_1577# 0.01595f
C1441 a_53376_2122# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C1442 a_26296_2002# pin 0.00146f
C1443 a_50912_2122# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1444 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_3.gated_control 0.17277f
C1445 a_15936_2122# swmatrix_Tgate_4.gated_control 0.01553f
C1446 a_38676_1577# enable 0.00577f
C1447 swmatrix_Tgate_0.gated_control a_40748_1577# 0
C1448 a_38636_2122# enable 0.00368f
C1449 a_13472_2122# swmatrix_Tgate_4.gated_control 0.01496f
C1450 a_40380_1580# ShiftReg_row_10_2$1_0.Q[7] 0.00101f
C1451 a_38776_2002# a_38676_1577# 0
C1452 a_37916_1580# a_38284_1577# 0.00194f
C1453 a_39912_1562# ShiftReg_row_10_2$1_0.Q[7] 0.00225f
C1454 a_44916_1577# pin 0
C1455 swmatrix_Tgate_3.gated_control vdd 1.84761f
C1456 a_38776_2002# a_38636_2122# 0.00109f
C1457 a_25804_1577# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1458 a_52860_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1459 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_1.gated_control 0.23535f
C1460 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1461 a_7232_2122# a_7476_1577# 0.01595f
C1462 a_18728_1562# pin 0
C1463 a_52392_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1464 a_24968_1562# a_26296_2002# 0.02403f
C1465 swmatrix_Tgate_7.gated_control a_25436_1580# 0
C1466 a_6716_1580# a_7576_2002# 0.00888f
C1467 a_40380_1580# vdd 0.42496f
C1468 a_7232_2122# a_7436_2122# 0.01151f
C1469 a_53228_1577# enable 0.0022f
C1470 a_39912_1562# vdd 1.0427f
C1471 ShiftReg_row_10_2$1_0.Q[8] a_51256_2002# 0.00242f
C1472 a_22176_2122# a_22028_2122# 0
C1473 a_21660_1580# a_22520_2002# 0.00888f
C1474 a_13676_2122# PHI_1 0.00534f
C1475 a_21192_1562# a_22520_2002# 0.02403f
C1476 swmatrix_Tgate_2.gated_control d_out 0.22358f
C1477 a_19712_2122# a_20056_2002# 0.57845f
C1478 a_21192_1562# a_19196_1580# 0
C1479 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_17401_1539# 0.0097f
C1480 a_1196_2122# enable 0.00368f
C1481 ShiftReg_row_10_2$1_0.Q[9] BUS[9] 0.01695f
C1482 a_34860_2122# swmatrix_Tgate_6.gated_control 0
C1483 a_59468_2122# vdd 0.00491f
C1484 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[3] 0
C1485 a_22520_2002# enable 0.0522f
C1486 a_57496_2002# vdd 0.32603f
C1487 a_19196_1580# enable 0.05108f
C1488 a_28760_2002# pin 0
C1489 ShiftReg_row_10_2$1_0.Q[6] PHI_1 0.05798f
C1490 a_57496_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1491 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C1492 a_25436_1580# pin 0
C1493 a_59860_1577# pin 0
C1494 a_3660_2122# vdd 0.01506f
C1495 swmatrix_Tgate_0.gated_control a_44524_1577# 0
C1496 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.08486f
C1497 a_41100_2122# enable 0.00368f
C1498 swmatrix_Tgate_0.gated_control a_41140_1577# 0
C1499 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1500 a_38284_2122# enable 0.00101f
C1501 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C1502 a_40896_2122# ShiftReg_row_10_2$1_0.Q[7] 0.11433f
C1503 a_43688_1562# BUS[8] 0.0057f
C1504 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C1505 a_9696_2122# a_9900_2122# 0.01151f
C1506 a_9180_1580# a_9548_2122# 0.00294f
C1507 a_49928_1562# vdd 1.00067f
C1508 a_26196_1577# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1509 a_7232_2122# a_7084_2122# 0
C1510 a_8712_1562# a_7576_2002# 0
C1511 a_57004_1577# enable 0.0022f
C1512 a_53376_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1513 a_53620_1577# enable 0.00579f
C1514 a_24968_1562# a_25436_1580# 0.30528f
C1515 a_40896_2122# vdd 0.55944f
C1516 a_38432_2122# vdd 0.56482f
C1517 a_22176_2122# a_22520_2002# 0.57845f
C1518 swmatrix_Tgate_5.gated_control enable 0.50846f
C1519 a_21192_1562# a_21660_1580# 0.30528f
C1520 a_16140_2122# PHI_1 0.00477f
C1521 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1522 ShiftReg_row_10_2$1_0.Q[2] a_13816_2002# 0.00242f
C1523 ShiftReg_row_10_2$1_0.Q[8] a_50396_1580# 0.36203f
C1524 a_13324_2122# PHI_1 0.00201f
C1525 a_19712_2122# a_19196_1580# 0.30053f
C1526 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C1527 a_50764_1577# BUS[9] 0
C1528 a_21660_1580# enable 0.05124f
C1529 a_21192_1562# enable 0.08694f
C1530 a_59960_2002# vdd 0.32887f
C1531 a_32536_2002# swmatrix_Tgate_6.gated_control 0.01121f
C1532 swmatrix_Tgate_6.gated_control pin 1.23291f
C1533 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[3] 0.01102f
C1534 a_56636_1580# vdd 0.42253f
C1535 a_27900_1580# pin 0.00113f
C1536 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_59960_2002# 0.00242f
C1537 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C1538 PHI_2 d_out 0.32019f
C1539 a_56636_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1540 a_27432_1562# pin 0.00138f
C1541 a_36121_1539# BUS[6] 0
C1542 a_3308_2122# vdd 0.00491f
C1543 a_40748_2122# enable 0.00101f
C1544 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42643f
C1545 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C1546 a_38776_2002# enable 0.05124f
C1547 a_41240_2002# a_41100_2122# 0.00109f
C1548 a_38432_2122# a_38284_1577# 0
C1549 a_31208_1562# swmatrix_Tgate_5.gated_control 0.00493f
C1550 a_45016_2002# pin 0.00146f
C1551 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C1552 a_37916_1580# a_38284_2122# 0.00294f
C1553 a_9696_2122# a_9548_2122# 0
C1554 a_9180_1580# a_10040_2002# 0.00888f
C1555 ShiftReg_row_10_2$1_0.Q[9] swmatrix_Tgate_1.gated_control 0.22418f
C1556 a_57396_1577# enable 0.00577f
C1557 a_8712_1562# a_10040_2002# 0.02403f
C1558 a_8712_1562# a_6716_1580# 0
C1559 a_57356_2122# enable 0.00368f
C1560 a_7232_2122# a_7576_2002# 0.57845f
C1561 pin BUS[9] 11.0719f
C1562 a_24968_1562# a_27432_1562# 0
C1563 a_992_2122# a_844_1577# 0
C1564 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C1565 swmatrix_Tgate_5.gated_control BUS[5] 0.86843f
C1566 a_46620_1580# a_46988_1577# 0.00194f
C1567 ShiftReg_row_10_2$1_0.Q[2] a_12956_1580# 0.36203f
C1568 a_47480_2002# a_47380_1577# 0
C1569 a_22176_2122# a_21660_1580# 0.30053f
C1570 a_31208_1562# enable 0.08752f
C1571 a_21192_1562# a_22176_2122# 0.07055f
C1572 a_15788_2122# PHI_1 0.00164f
C1573 a_19712_2122# a_21192_1562# 0.00268f
C1574 a_13816_2002# PHI_1 0.01314f
C1575 a_51156_1577# BUS[9] 0
C1576 a_37448_1562# pin 0
C1577 a_35000_2002# swmatrix_Tgate_6.gated_control 0.01014f
C1578 a_22176_2122# enable 0.11443f
C1579 a_31676_1580# swmatrix_Tgate_6.gated_control 0.00804f
C1580 a_59100_1580# vdd 0.42496f
C1581 a_19712_2122# enable 0.11055f
C1582 a_51116_2122# BUS[9] 0
C1583 a_58632_1562# vdd 1.0427f
C1584 enable BUS[5] 0.2115f
C1585 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_59100_1580# 0.36162f
C1586 a_28416_2122# pin 0.00251f
C1587 a_58632_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1588 a_4921_1539# pin 0
C1589 a_25952_2122# pin 0.00138f
C1590 a_32396_2122# PHI_1 0.00534f
C1591 a_34508_1577# BUS[6] 0
C1592 a_3800_2002# vdd 0.32879f
C1593 a_41240_2002# enable 0.0522f
C1594 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1595 a_2472_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1596 a_37916_1580# enable 0.05108f
C1597 vdd BUS[6] 0.56053f
C1598 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1599 ShiftReg_row_10_2$1_0.Q[9] PHI_1 0.05798f
C1600 a_38432_2122# a_38676_1577# 0.01595f
C1601 a_47480_2002# pin 0
C1602 a_44156_1580# pin 0
C1603 a_38432_2122# a_38636_2122# 0.01151f
C1604 a_37916_1580# a_38776_2002# 0.00888f
C1605 a_9696_2122# a_10040_2002# 0.57845f
C1606 ShiftReg_row_10_2$1_0.Q[9] a_56168_1562# 0.16779f
C1607 a_59820_2122# enable 0.00368f
C1608 a_26296_2002# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1609 a_8712_1562# a_9180_1580# 0.30528f
C1610 a_50764_1577# swmatrix_Tgate_1.gated_control 0
C1611 a_7232_2122# a_6716_1580# 0.30053f
C1612 a_57004_2122# enable 0.00101f
C1613 a_24968_1562# a_25952_2122# 0.07055f
C1614 a_17401_1539# PHI_2 0
C1615 a_992_2122# a_1236_1577# 0.01595f
C1616 a_12488_1562# BUS[3] 0.0057f
C1617 a_10040_2002# a_9940_1577# 0
C1618 swmatrix_Tgate_6.gated_control swmatrix_Tgate_0.gated_control 0.01259f
C1619 ShiftReg_row_10_2$1_0.Q[8] a_50912_2122# 0.01552f
C1620 PHI_2 BUS[3] 0.11252f
C1621 a_47136_2122# a_46988_1577# 0
C1622 a_9180_1580# a_9548_1577# 0.00194f
C1623 a_16280_2002# PHI_1 0.01261f
C1624 a_6248_1562# BUS[2] 0.0057f
C1625 a_12956_1580# PHI_1 0.0533f
C1626 a_53580_2122# BUS[9] 0.00104f
C1627 a_34140_1580# swmatrix_Tgate_6.gated_control 0.00668f
C1628 a_43688_1562# swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1629 a_33672_1562# swmatrix_Tgate_6.gated_control 0.00985f
C1630 a_50764_2122# BUS[9] 0
C1631 a_59616_2122# vdd 0.55944f
C1632 a_57152_2122# vdd 0.56482f
C1633 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_59616_2122# 0.01536f
C1634 ShiftReg_row_10_2$1_0.Q[2] pin 0.01491f
C1635 swmatrix_Tgate_3.gated_control enable 0.50846f
C1636 ShiftReg_row_10_2$1_0.Q[5] ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1637 a_57152_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C1638 a_3308_1577# pin 0
C1639 a_34860_2122# PHI_1 0.00477f
C1640 a_34900_1577# BUS[6] 0
C1641 a_32044_2122# PHI_1 0.00201f
C1642 a_2940_1580# vdd 0.42489f
C1643 a_2472_1562# a_3800_2002# 0.02403f
C1644 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C1645 a_57004_1577# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1646 swmatrix_Tgate_1.gated_control pin 1.23291f
C1647 ShiftReg_row_10_2$1_0.Q[4] ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C1648 a_40380_1580# enable 0.05124f
C1649 a_39912_1562# enable 0.08694f
C1650 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_22028_1577# 0
C1651 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1652 a_40380_1580# a_40748_2122# 0.00294f
C1653 a_40896_2122# a_41100_2122# 0.01151f
C1654 a_46620_1580# pin 0.00113f
C1655 a_9696_2122# a_9180_1580# 0.30053f
C1656 a_46152_1562# pin 0.00138f
C1657 a_38432_2122# a_38284_2122# 0
C1658 a_39912_1562# a_38776_2002# 0
C1659 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_3800_2002# 0.00242f
C1660 a_28760_2002# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C1661 a_8712_1562# a_9696_2122# 0.07055f
C1662 a_51156_1577# swmatrix_Tgate_1.gated_control 0
C1663 a_7232_2122# a_8712_1562# 0.00268f
C1664 ShiftReg_row_10_2$1_0.Q[4] PHI_2 0.63578f
C1665 a_25436_1580# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1666 a_51116_2122# swmatrix_Tgate_1.gated_control 0
C1667 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.08552f
C1668 a_59468_2122# enable 0.00101f
C1669 a_57496_2002# enable 0.05124f
C1670 swmatrix_Tgate_7.gated_control PHI_1 0.01086f
C1671 a_15788_1577# PHI_2 0
C1672 ShiftReg_row_10_2$1_0.Q[2] a_13472_2122# 0.01552f
C1673 a_9696_2122# a_9548_1577# 0
C1674 a_15420_1580# PHI_1 0.01277f
C1675 a_37448_1562# swmatrix_Tgate_0.gated_control 0.01486f
C1676 a_47136_2122# a_47380_1577# 0.01595f
C1677 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C1678 a_14952_1562# PHI_1 0.01733f
C1679 a_3660_2122# enable 0.00368f
C1680 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C1681 ShiftReg_row_10_2$1_0.Q[1] vdd 0.57762f
C1682 a_8_1562# PHI_2 0.02723f
C1683 a_34656_2122# swmatrix_Tgate_6.gated_control 0.01553f
C1684 swmatrix_Tgate_4.gated_control BUS[2] 0.00566f
C1685 a_53228_2122# BUS[9] 0
C1686 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C1687 a_51256_2002# BUS[9] 0.0117f
C1688 a_32192_2122# swmatrix_Tgate_6.gated_control 0.01496f
C1689 a_59100_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1690 a_49928_1562# enable 0.08752f
C1691 a_34508_2122# PHI_1 0.00164f
C1692 a_56636_1580# a_57004_1577# 0.00194f
C1693 a_58632_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1694 a_57496_2002# a_57396_1577# 0
C1695 PHI_1 pin 0.0015f
C1696 a_3700_1577# pin 0
C1697 a_57496_2002# a_57356_2122# 0.00109f
C1698 a_992_2122# pin 0.00343f
C1699 a_32536_2002# PHI_1 0.01314f
C1700 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[7] 0.10774f
C1701 a_3456_2122# vdd 0.56033f
C1702 a_2472_1562# a_2940_1580# 0.30528f
C1703 ShiftReg_row_10_2$1_0.Q[4] a_23641_1539# 0.00241f
C1704 a_43688_1562# a_45016_2002# 0.02403f
C1705 a_56168_1562# pin 0
C1706 swmatrix_Tgate_0.gated_control a_44156_1580# 0
C1707 a_57396_1577# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1708 a_40896_2122# enable 0.11443f
C1709 a_38432_2122# enable 0.11055f
C1710 swmatrix_Tgate_6.gated_control swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C1711 a_40896_2122# a_40748_2122# 0
C1712 a_40380_1580# a_41240_2002# 0.00888f
C1713 a_47136_2122# pin 0.00251f
C1714 a_39912_1562# a_41240_2002# 0.02403f
C1715 a_3308_1577# BUS[1] 0
C1716 a_39912_1562# a_37916_1580# 0
C1717 a_51116_2122# PHI_1 0.00534f
C1718 a_38432_2122# a_38776_2002# 0.57845f
C1719 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_36121_1539# 0.0097f
C1720 a_44672_2122# pin 0.00138f
C1721 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_2940_1580# 0.36162f
C1722 a_27900_1580# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C1723 a_53580_2122# swmatrix_Tgate_1.gated_control 0
C1724 a_27432_1562# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C1725 a_59960_2002# enable 0.0522f
C1726 a_19564_1577# PHI_2 0
C1727 a_56636_1580# enable 0.05108f
C1728 a_16180_1577# PHI_2 0
C1729 a_24968_1562# PHI_1 0.70141f
C1730 a_9696_2122# a_9940_1577# 0.01595f
C1731 a_15936_2122# PHI_1 0.01804f
C1732 a_3308_2122# enable 0.00101f
C1733 a_13472_2122# PHI_1 0.01882f
C1734 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1735 swmatrix_Tgate_2.gated_control vdd 1.85047f
C1736 a_53720_2002# BUS[9] 0.01161f
C1737 a_2472_1562# ShiftReg_row_10_2$1_0.Q[1] 0.00225f
C1738 a_50396_1580# BUS[9] 0.00688f
C1739 a_36121_1539# PHI_2 0
C1740 a_1336_2002# a_1236_1577# 0
C1741 a_13816_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1742 a_59616_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1743 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_2.gated_control 0.23535f
C1744 a_7476_1577# pin 0
C1745 swmatrix_Tgate_8.gated_control vdd 1.84484f
C1746 a_35000_2002# PHI_1 0.01261f
C1747 a_31676_1580# PHI_1 0.0533f
C1748 a_2472_1562# a_3456_2122# 0.07055f
C1749 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[1] 0.01102f
C1750 a_43688_1562# a_44156_1580# 0.30528f
C1751 a_40896_2122# a_41240_2002# 0.57845f
C1752 a_39912_1562# a_40380_1580# 0.30528f
C1753 a_3700_1577# BUS[1] 0
C1754 a_53580_2122# PHI_1 0.00477f
C1755 a_992_2122# BUS[1] 0.01972f
C1756 a_50764_2122# PHI_1 0.00201f
C1757 PHI_1 BUS[1] 0.09541f
C1758 a_38432_2122# a_37916_1580# 0.30053f
C1759 a_28416_2122# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C1760 a_25952_2122# swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1761 a_59100_1580# enable 0.05124f
C1762 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_3456_2122# 0.01536f
C1763 a_58632_1562# enable 0.08694f
C1764 a_19956_1577# PHI_2 0
C1765 pin BUS[10] 11.0719f
C1766 a_51256_2002# swmatrix_Tgate_1.gated_control 0.01121f
C1767 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[6] 0.01102f
C1768 a_19916_2122# PHI_2 0.00411f
C1769 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1770 a_3800_2002# enable 0.0522f
C1771 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C1772 a_61081_1539# d_out 0.00241f
C1773 a_8_1562# D_in 0.15891f
C1774 swmatrix_Tgate_0.gated_control PHI_1 0.01086f
C1775 ShiftReg_row_10_2$1_0.Q[7] PHI_2 0.63578f
C1776 a_52860_1580# BUS[9] 0.01336f
C1777 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_16280_2002# 0.00242f
C1778 a_34508_1577# PHI_2 0
C1779 a_12956_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C1780 a_52392_1562# BUS[9] 0.02637f
C1781 a_59960_2002# a_59820_2122# 0.00109f
C1782 enable BUS[6] 0.2115f
C1783 a_57152_2122# a_57004_1577# 0
C1784 a_49928_1562# swmatrix_Tgate_3.gated_control 0.00493f
C1785 a_34140_1580# PHI_1 0.01277f
C1786 ShiftReg_row_10_2$1_0.Q[7] BUS[7] 0.01695f
C1787 a_12488_1562# vdd 1.00067f
C1788 a_56636_1580# a_57004_2122# 0.00294f
C1789 vdd PHI_2 4.67187f
C1790 a_33672_1562# PHI_1 0.01733f
C1791 a_476_1580# PHI_2 0.03321f
C1792 ShiftReg_row_10_2$1_0.Q[4] a_25804_1577# 0
C1793 a_43688_1562# a_46152_1562# 0
C1794 a_57496_2002# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1795 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C1796 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[2] 0.10774f
C1797 a_40896_2122# a_40380_1580# 0.30053f
C1798 vdd BUS[7] 0.56053f
C1799 a_53228_2122# PHI_1 0.00164f
C1800 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C1801 a_39912_1562# a_40896_2122# 0.07055f
C1802 a_1336_2002# pin 0
C1803 a_38432_2122# a_39912_1562# 0.00268f
C1804 a_51256_2002# PHI_1 0.01314f
C1805 a_53720_2002# swmatrix_Tgate_1.gated_control 0.01014f
C1806 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C1807 a_50396_1580# swmatrix_Tgate_1.gated_control 0.00804f
C1808 a_22380_2122# PHI_2 0.00422f
C1809 a_59616_2122# enable 0.11443f
C1810 a_57152_2122# enable 0.11055f
C1811 a_19564_2122# PHI_2 0
C1812 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_7.gated_control 0.33472f
C1813 a_31208_1562# BUS[6] 0.0057f
C1814 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1815 PHI_2 BUS[4] 0.11252f
C1816 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00204f
C1817 a_844_2122# BUS[1] 0
C1818 a_2940_1580# enable 0.05124f
C1819 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1820 a_53376_2122# BUS[9] 0.01571f
C1821 a_38284_1577# PHI_2 0
C1822 a_50912_2122# BUS[9] 0.0191f
C1823 a_43688_1562# PHI_1 0.70141f
C1824 a_8_1562# swmatrix_Tgate_9.gated_control 0.01276f
C1825 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_15420_1580# 0.36162f
C1826 a_34900_1577# PHI_2 0
C1827 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1828 a_14952_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C1829 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_2.gated_control 0.33472f
C1830 a_34656_2122# PHI_1 0.01804f
C1831 a_57152_2122# a_57396_1577# 0.01595f
C1832 a_7576_2002# pin 0.00146f
C1833 a_32192_2122# PHI_1 0.01882f
C1834 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C1835 a_56636_1580# a_57496_2002# 0.00888f
C1836 a_38284_1577# BUS[7] 0
C1837 a_57152_2122# a_57356_2122# 0.01151f
C1838 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C1839 a_2472_1562# PHI_2 0.60119f
C1840 a_54841_1539# PHI_2 0
C1841 a_59960_2002# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C1842 a_43688_1562# a_44672_2122# 0.07055f
C1843 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C1844 a_56636_1580# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1845 a_53720_2002# PHI_1 0.01261f
C1846 a_23641_1539# BUS[4] 0
C1847 a_50396_1580# PHI_1 0.0533f
C1848 a_52860_1580# swmatrix_Tgate_1.gated_control 0.00668f
C1849 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_2 0.45413f
C1850 ShiftReg_row_10_2$1_0.Q[1] enable 0.513f
C1851 a_8_1562# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1852 a_22028_2122# PHI_2 0
C1853 a_52392_1562# swmatrix_Tgate_1.gated_control 0.00985f
C1854 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C1855 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_24968_1562# 0
C1856 a_20056_2002# PHI_2 0.03207f
C1857 a_1336_2002# BUS[1] 0.01428f
C1858 swmatrix_Tgate_4.gated_control a_17401_1539# 0.00113f
C1859 a_18728_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C1860 ShiftReg_row_10_2$1_0.Q[8] ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C1861 a_3456_2122# enable 0.11443f
C1862 ShiftReg_row_10_2$1_0.Q[5] vdd 0.57779f
C1863 swmatrix_Tgate_4.gated_control BUS[3] 0.86843f
C1864 ShiftReg_row_10_2$1_0.Q[7] ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.01068f
C1865 a_38676_1577# PHI_2 0
C1866 a_16280_2002# ShiftReg_row_10_2$1_0.Q[3] 0.25874f
C1867 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_40748_1577# 0
C1868 a_38636_2122# PHI_2 0.00411f
C1869 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[8] 0
C1870 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_15936_2122# 0.01536f
C1871 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vdd 0.42852f
C1872 a_13472_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C1873 a_57004_1577# swmatrix_Tgate_2.gated_control 0
C1874 a_10040_2002# pin 0
C1875 a_59616_2122# a_59820_2122# 0.01151f
C1876 a_59100_1580# a_59468_2122# 0.00294f
C1877 a_38676_1577# BUS[7] 0
C1878 a_6716_1580# pin 0
C1879 a_38636_2122# BUS[7] 0
C1880 a_58632_1562# a_57496_2002# 0
C1881 a_57152_2122# a_57004_2122# 0
C1882 vdd D_in 0.18311f
C1883 a_476_1580# D_in 0.36155f
C1884 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C1885 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C1886 swmatrix_Tgate_0.gated_control swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C1887 a_53228_1577# PHI_2 0
C1888 a_59100_1580# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C1889 a_58632_1562# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00397f
C1890 ShiftReg_row_10_2$1_0.Q[2] BUS[2] 0.01695f
C1891 a_22028_1577# BUS[4] 0
C1892 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_8.gated_control 0.33472f
C1893 a_52860_1580# PHI_1 0.01277f
C1894 a_52392_1562# PHI_1 0.01733f
C1895 a_1196_2122# PHI_2 0.00411f
C1896 swmatrix_Tgate_2.gated_control enable 0.50433f
C1897 a_3800_2002# a_3660_2122# 0.00109f
C1898 a_53376_2122# swmatrix_Tgate_1.gated_control 0.01553f
C1899 a_22520_2002# PHI_2 0.03174f
C1900 a_50912_2122# swmatrix_Tgate_1.gated_control 0.01496f
C1901 a_19196_1580# PHI_2 0.03321f
C1902 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00347f
C1903 ShiftReg_row_10_2$1_0.Q[3] swmatrix_Tgate_7.gated_control 0.17277f
C1904 swmatrix_Tgate_8.gated_control enable 0.50846f
C1905 swmatrix_Tgate_4.gated_control a_15788_1577# 0
C1906 a_15420_1580# ShiftReg_row_10_2$1_0.Q[3] 0.00101f
C1907 a_41100_2122# PHI_2 0.00422f
C1908 ShiftReg_row_10_2$1_0.Q[7] a_42361_1539# 0.00241f
C1909 a_57396_1577# swmatrix_Tgate_2.gated_control 0
C1910 a_14952_1562# ShiftReg_row_10_2$1_0.Q[3] 0.00225f
C1911 a_13816_2002# a_13716_1577# 0
C1912 a_12956_1580# a_13324_1577# 0.00194f
C1913 a_38284_2122# PHI_2 0
C1914 a_13816_2002# a_13676_2122# 0.00109f
C1915 a_59100_1580# a_59960_2002# 0.00888f
C1916 a_57356_2122# swmatrix_Tgate_2.gated_control 0
C1917 a_59616_2122# a_59468_2122# 0
C1918 a_58632_1562# a_59960_2002# 0.02403f
C1919 a_9180_1580# pin 0.00113f
C1920 a_41100_2122# BUS[7] 0.00104f
C1921 a_27900_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1922 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_5.gated_control 0.23535f
C1923 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_54841_1539# 0.0097f
C1924 a_57152_2122# a_57496_2002# 0.57845f
C1925 a_58632_1562# a_56636_1580# 0
C1926 a_8712_1562# pin 0.00138f
C1927 a_27432_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1928 a_38284_2122# BUS[7] 0
C1929 swmatrix_Tgate_9.gated_control vdd 1.83165f
C1930 a_57004_1577# PHI_2 0
C1931 a_476_1580# swmatrix_Tgate_9.gated_control 0.00784f
C1932 ShiftReg_row_10_2$1_0.Q[3] pin 0.01491f
C1933 a_59616_2122# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00475f
C1934 ShiftReg_row_10_2$1_0.Q[4] a_26296_2002# 0.00242f
C1935 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C1936 a_53620_1577# PHI_2 0
C1937 a_7084_1577# BUS[2] 0
C1938 a_57152_2122# swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1939 a_18728_1562# swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1940 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_12488_1562# 0
C1941 a_22420_1577# BUS[4] 0
C1942 a_53376_2122# PHI_1 0.01804f
C1943 swmatrix_Tgate_5.gated_control PHI_2 0.31095f
C1944 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C1945 PHI_1 BUS[2] 0.09486f
C1946 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN pin 0
C1947 a_12488_1562# swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1948 a_50912_2122# PHI_1 0.01882f
C1949 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C1950 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q D_in 0.01068f
C1951 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C1952 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C1953 a_21660_1580# PHI_2 0.07395f
C1954 a_32536_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C1955 a_21192_1562# PHI_2 0.60119f
C1956 a_32044_1577# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1957 swmatrix_Tgate_4.gated_control a_19564_1577# 0
C1958 a_12488_1562# enable 0.08752f
C1959 swmatrix_Tgate_4.gated_control a_16180_1577# 0
C1960 PHI_2 enable 1.35356f
C1961 a_26156_2122# vdd 0.01506f
C1962 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.08448f
C1963 a_476_1580# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1964 a_15936_2122# ShiftReg_row_10_2$1_0.Q[3] 0.11433f
C1965 a_40748_2122# PHI_2 0
C1966 a_38776_2002# PHI_2 0.03207f
C1967 a_59820_2122# swmatrix_Tgate_2.gated_control 0
C1968 enable BUS[7] 0.2115f
C1969 a_59616_2122# a_59960_2002# 0.57845f
C1970 a_9696_2122# pin 0.00251f
C1971 a_58632_1562# a_59100_1580# 0.30528f
C1972 a_28416_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C1973 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09546f
C1974 a_7232_2122# pin 0.00138f
C1975 ShiftReg_row_10_2$1_0.Q[8] vdd 0.57779f
C1976 a_40748_2122# BUS[7] 0
C1977 a_57152_2122# a_56636_1580# 0.30053f
C1978 a_38776_2002# BUS[7] 0.0117f
C1979 a_6248_1562# vdd 1.00067f
C1980 a_2472_1562# swmatrix_Tgate_9.gated_control 0.00985f
C1981 a_57396_1577# PHI_2 0
C1982 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q ShiftReg_row_10_2$1_0.Q[9] 0.01102f
C1983 ShiftReg_row_10_2$1_0.Q[4] a_25436_1580# 0.36203f
C1984 a_9940_1577# pin 0
C1985 a_57356_2122# PHI_2 0.00411f
C1986 a_7476_1577# BUS[2] 0
C1987 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q BUS[5] 0.10774f
C1988 vdd BUS[8] 0.56053f
C1989 a_7436_2122# BUS[2] 0
C1990 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C1991 a_31208_1562# PHI_2 0.02762f
C1992 a_23641_1539# enable 0.00398f
C1993 a_2940_1580# a_3308_2122# 0.00294f
C1994 a_3456_2122# a_3660_2122# 0.01151f
C1995 a_22176_2122# PHI_2 0.04011f
C1996 a_2940_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C1997 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_35000_2002# 0.00242f
C1998 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_9.gated_control 0.23535f
C1999 a_19712_2122# PHI_2 0.04895f
C2000 a_31676_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0
C2001 PHI_2 BUS[5] 0.11252f
C2002 a_32436_1577# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2003 a_28620_2122# vdd 0.01506f
C2004 a_25804_2122# vdd 0.00491f
C2005 ShiftReg_row_10_2$1_0.Q[7] a_44524_1577# 0
C2006 a_16280_2002# a_16140_2122# 0.00109f
C2007 a_41240_2002# PHI_2 0.03174f
C2008 a_2472_1562# swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00368f
C2009 a_37916_1580# PHI_2 0.03321f
C2010 a_13472_2122# a_13324_1577# 0
C2011 a_12956_1580# a_13324_2122# 0.00294f
C2012 a_59616_2122# a_59100_1580# 0.30053f
C2013 a_57496_2002# swmatrix_Tgate_2.gated_control 0.01121f
C2014 a_58632_1562# a_59616_2122# 0.07055f
C2015 ShiftReg_row_10_2$1_0.Q[5] swmatrix_Tgate_5.gated_control 0.22418f
C2016 a_41240_2002# BUS[7] 0.01161f
C2017 a_57152_2122# a_58632_1562# 0.00268f
C2018 a_37916_1580# BUS[7] 0.00688f
C2019 swmatrix_Tgate_2.gated_control swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C2020 a_59820_2122# PHI_2 0.00422f
C2021 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00188f
C2022 a_22520_2002# a_22420_1577# 0
C2023 a_57004_2122# PHI_2 0
C2024 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN swmatrix_Tgate_0.gated_control 0.33472f
C2025 a_21660_1580# a_22028_1577# 0.00194f
C2026 a_13716_1577# pin 0
C2027 swmatrix_Tgate_4.gated_control vdd 1.84761f
C2028 ShiftReg_row_10_2$1_0.Q[1] ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.08575f
C2029 a_9900_2122# BUS[2] 0.00104f
C2030 ShiftReg_row_10_2$1_0.Q[5] enable 0.513f
C2031 a_7084_2122# BUS[2] 0
C2032 a_22028_1577# enable 0.0022f
C2033 a_3456_2122# a_3308_2122# 0
C2034 a_2940_1580# a_3800_2002# 0.00888f
C2035 a_1196_2122# swmatrix_Tgate_9.gated_control 0
C2036 a_3456_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0.00144f
C2037 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_34140_1580# 0.36162f
C2038 ShiftReg_row_10_2$1_0.Q[6] pin 0.01491f
C2039 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN enable 0.65271f
C2040 a_33672_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.16689f
C2041 D_in enable 0.13355f
C2042 swmatrix_Tgate_3.gated_control PHI_2 0.31095f
C2043 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q enable 0.20415f
C2044 PHI_1 d_out 0.03331f
C2045 a_28268_2122# vdd 0.00491f
C2046 a_26296_2002# vdd 0.32603f
C2047 a_40380_1580# PHI_2 0.07395f
C2048 a_13472_2122# a_13716_1577# 0.01595f
C2049 swmatrix_Tgate_3.gated_control BUS[7] 0.00566f
C2050 a_39912_1562# PHI_2 0.60119f
C2051 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q pin 0
C2052 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_59468_1577# 0
C2053 a_59960_2002# swmatrix_Tgate_2.gated_control 0.01014f
C2054 a_12956_1580# a_13816_2002# 0.00888f
C2055 a_13472_2122# a_13676_2122# 0.01151f
C2056 ShiftReg_row_10_2$1_0.Q[5] a_31208_1562# 0.16779f
C2057 a_25804_1577# swmatrix_Tgate_5.gated_control 0
C2058 a_56636_1580# swmatrix_Tgate_2.gated_control 0.00804f
C2059 a_40380_1580# BUS[7] 0.01336f
C2060 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C2061 a_39912_1562# BUS[7] 0.02637f
C2062 a_44876_2122# vdd 0.01506f
C2063 a_59468_2122# PHI_2 0
C2064 a_3800_2002# ShiftReg_row_10_2$1_0.Q[1] 0.25874f
C2065 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_43688_1562# 0
C2066 a_22176_2122# a_22028_1577# 0
C2067 a_57496_2002# PHI_2 0.03207f
C2068 ShiftReg_row_10_2$1_0.Q[4] a_25952_2122# 0.01552f
C2069 ShiftReg_row_10_2$1_0.Q[5] BUS[5] 0.01695f
C2070 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C2071 a_18728_1562# vdd 1.00067f
C2072 a_9548_2122# BUS[2] 0
C2073 swmatrix_Tgate_6.gated_control a_36121_1539# 0.00113f
C2074 a_37448_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.00116f
C2075 a_7576_2002# BUS[2] 0.0117f
C2076 a_25804_1577# enable 0.0022f
C2077 a_3660_2122# PHI_2 0.00422f
C2078 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_2 0.00169f
C2079 a_22420_1577# enable 0.00579f
C2080 a_3456_2122# a_3800_2002# 0.57845f
C2081 a_35000_2002# ShiftReg_row_10_2$1_0.Q[6] 0.25874f
C2082 ShiftReg_row_10_2$1_0.Q[7] swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2083 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q a_34656_2122# 0.01536f
C2084 a_32192_2122# ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.09501f
C2085 a_28660_1577# pin 0
C2086 a_32536_2002# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2087 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN pin 1.57433f
C2088 a_49928_1562# PHI_2 0.02762f
C2089 a_42361_1539# enable 0.00398f
C2090 a_28760_2002# vdd 0.32887f
C2091 swmatrix_Tgate_9.gated_control enable 0.51127f
C2092 a_25436_1580# vdd 0.42253f
C2093 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vdd 5.086f
C2094 a_18728_1562# BUS[4] 0.0057f
C2095 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN a_61081_1539# 0.0097f
C2096 a_40896_2122# PHI_2 0.04011f
C2097 a_15420_1580# a_15788_2122# 0.00294f
C2098 a_15936_2122# a_16140_2122# 0.01151f
C2099 a_59100_1580# swmatrix_Tgate_2.gated_control 0.00668f
C2100 a_38432_2122# PHI_2 0.04895f
C2101 a_14952_1562# a_13816_2002# 0
C2102 a_58632_1562# swmatrix_Tgate_2.gated_control 0.00985f
C2103 a_13472_2122# a_13324_2122# 0
C2104 a_26196_1577# swmatrix_Tgate_5.gated_control 0
C2105 a_40896_2122# BUS[7] 0.01571f
C2106 a_49928_1562# swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2107 a_47340_2122# vdd 0.01506f
C2108 a_26156_2122# swmatrix_Tgate_5.gated_control 0
C2109 a_44524_2122# vdd 0.00491f
C2110 a_38432_2122# BUS[7] 0.0191f
C2111 a_2940_1580# ShiftReg_row_10_2$1_0.Q[1] 0.00101f
C2112 d_out BUS[10] 0.01695f
C2113 a_59960_2002# PHI_2 0.03174f
C2114 a_22176_2122# a_22420_1577# 0.01595f
C2115 a_56636_1580# PHI_2 0.03321f
C2116 a_13816_2002# pin 0.00146f
C2117 a_10040_2002# BUS[2] 0.01161f
C2118 a_25804_1577# BUS[5] 0
C2119 ShiftReg_row_10_2$1_0.Q[6] swmatrix_Tgate_0.gated_control 0.17277f
C2120 a_6716_1580# BUS[2] 0.00688f
C2121 PHI_1 BUS[3] 0.09486f
C2122 a_26196_1577# enable 0.00577f
C2123 swmatrix_Tgate_6.gated_control a_34508_1577# 0
C2124 a_3456_2122# a_2940_1580# 0.30053f
C2125 a_26156_2122# enable 0.00368f
C2126 a_3308_2122# PHI_2 0
C2127 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN enable 0.09559f
C2128 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_2 0.03773f
C2129 a_32436_1577# pin 0
C2130 a_34140_1580# ShiftReg_row_10_2$1_0.Q[6] 0.00101f
C2131 a_33672_1562# ShiftReg_row_10_2$1_0.Q[6] 0.00225f
C2132 a_32536_2002# a_32436_1577# 0
C2133 a_31676_1580# a_32044_1577# 0.00194f
C2134 a_11161_1539# BUS[2] 0
C2135 ShiftReg_row_10_2$1_0.Q[1] swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2136 swmatrix_Tgate_6.gated_control vdd 1.84761f
C2137 a_32536_2002# a_32396_2122# 0.00109f
C2138 a_35000_2002# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.0016f
C2139 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q swmatrix_Tgate_3.gated_control 0.23535f
C2140 ShiftReg_row_10_2$1_0.Q[8] enable 0.513f
C2141 a_46620_1580# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C2142 a_31676_1580# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0
C2143 a_27900_1580# vdd 0.42496f
C2144 a_46152_1562# ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN 0
C2145 a_40748_1577# enable 0.0022f
C2146 swmatrix_Tgate_4.gated_control a_19196_1580# 0
C2147 a_18728_1562# a_20056_2002# 0.02403f
C2148 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vdd 0.34474f
C2149 a_27432_1562# vdd 1.0427f
C2150 a_6248_1562# enable 0.08752f
C2151 a_15420_1580# a_16280_2002# 0.00888f
C2152 ShiftReg_row_10_2$1_0.Q[9] pin 0.01491f
C2153 a_15936_2122# a_15788_2122# 0
C2154 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN PHI_1 0
C2155 a_14952_1562# a_16280_2002# 0.02403f
C2156 enable BUS[8] 0.2115f
C2157 ShiftReg_row_10_2$1_0.Q[7] a_45016_2002# 0.00242f
C2158 a_13472_2122# a_13816_2002# 0.57845f
C2159 a_59616_2122# swmatrix_Tgate_2.gated_control 0.01553f
C2160 a_14952_1562# a_12956_1580# 0
C2161 a_57152_2122# swmatrix_Tgate_2.gated_control 0.01496f
C2162 a_28620_2122# swmatrix_Tgate_5.gated_control 0
C2163 a_1236_1577# pin 0
C2164 a_46988_2122# vdd 0.00491f
C2165 a_45016_2002# vdd 0.32603f
C2166 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN BUS[6] 0
C2167 a_3456_2122# ShiftReg_row_10_2$1_0.Q[1] 0.11433f
C2168 ShiftReg_row_10_2$1_0.Q[4] PHI_1 0.05798f
C2169 a_59100_1580# PHI_2 0.07395f
C2170 a_16280_2002# pin 0
C2171 vdd BUS[9] 0.56053f
C2172 a_58632_1562# PHI_2 0.60119f
C2173 a_12956_1580# pin 0
C2174 a_26196_1577# BUS[5] 0
C2175 a_51256_2002# ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q 0.2556f
C2176 a_26156_2122# BUS[5] 0
C2177 a_9180_1580# BUS[2] 0.01336f
C2178 a_8712_1562# BUS[2] 0.02637f
C2179 swmatrix_Tgate_6.gated_control a_38284_1577# 0
C2180 a_28620_2122# enable 0.00368f
C2181 swmatrix_Tgate_6.gated_control a_34900_1577# 0
C2182 a_25804_2122# enable 0.00101f
C2183 a_844_1577# BUS[1] 0
C2184 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN PHI_1 0.02073f
C2185 a_3800_2002# PHI_2 0.03174f
C2186 a_61081_1539# enable 0.00398f
C2187 a_34656_2122# ShiftReg_row_10_2$1_0.Q[6] 0.11433f
C2188 swmatrix_Tgate_0.gated_control swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00518f
C2189 a_8_1562# PHI_1 0.70141f
C2190 a_8_1562# a_992_2122# 0.07055f
C2191 a_9548_1577# BUS[2] 0
C2192 a_37448_1562# vdd 1.00067f
C2193 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q PHI_1 0.01369f
C2194 PHI_2 BUS[6] 0.11252f
C2195 swmatrix_Tgate_4.gated_control swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.88137f
C2196 a_44524_1577# enable 0.0022f
C2197 a_34140_1580# swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN 0.00147f
C2198 BUS[10] vss 3.8004f
C2199 BUS[9] vss 3.79505f
C2200 BUS[8] vss 3.79505f
C2201 BUS[7] vss 3.79505f
C2202 BUS[6] vss 3.79505f
C2203 BUS[5] vss 3.79505f
C2204 BUS[4] vss 3.79505f
C2205 BUS[3] vss 3.79505f
C2206 BUS[2] vss 3.79505f
C2207 BUS[1] vss 4.14151f
C2208 pin vss 27.07676f
C2209 d_out vss 0.97418f
C2210 enable vss 24.46754f
C2211 PHI_2 vss 19.5562f
C2212 D_in vss 0.47925f
C2213 PHI_1 vss 29.7212f
C2214 vdd vss 0.29571p
C2215 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84863f
C2216 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2217 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2218 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2219 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2220 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2221 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2222 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84749f
C2223 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.84796f
C2224 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN vss 1.85974f
C2225 a_61081_1539# vss 0.0072f
C2226 a_59468_1577# vss 0.0042f
C2227 a_59860_1577# vss 0.0095f
C2228 swmatrix_Tgate_2.gated_control vss 3.21482f
C2229 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.77555f
C2230 a_57004_1577# vss 0.0042f
C2231 a_57396_1577# vss 0.0095f
C2232 a_59960_2002# vss 0.41829f
C2233 a_59100_1580# vss 0.52799f
C2234 a_59616_2122# vss 1.12757f
C2235 ShiftReg_row_10_2$1_0.DFF_2phase_1_0.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2236 a_54841_1539# vss 0.0072f
C2237 a_53228_1577# vss 0.0042f
C2238 a_53620_1577# vss 0.0095f
C2239 a_57496_2002# vss 0.42109f
C2240 a_56636_1580# vss 0.53063f
C2241 a_58632_1562# vss 1.18067f
C2242 a_57152_2122# vss 1.14287f
C2243 swmatrix_Tgate_1.gated_control vss 3.1994f
C2244 a_56168_1562# vss 1.1833f
C2245 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2246 ShiftReg_row_10_2$1_0.Q[9] vss 1.42957f
C2247 a_50764_1577# vss 0.0042f
C2248 a_51156_1577# vss 0.0095f
C2249 a_53720_2002# vss 0.41829f
C2250 a_52860_1580# vss 0.52799f
C2251 a_53376_2122# vss 1.12757f
C2252 ShiftReg_row_10_2$1_0.DFF_2phase_1_1.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2253 a_48601_1539# vss 0.0072f
C2254 a_46988_1577# vss 0.0042f
C2255 a_47380_1577# vss 0.0095f
C2256 a_51256_2002# vss 0.42109f
C2257 a_50396_1580# vss 0.53063f
C2258 a_52392_1562# vss 1.18067f
C2259 a_50912_2122# vss 1.14287f
C2260 swmatrix_Tgate_3.gated_control vss 3.1994f
C2261 a_49928_1562# vss 1.1833f
C2262 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2263 ShiftReg_row_10_2$1_0.Q[8] vss 1.42957f
C2264 a_44524_1577# vss 0.0042f
C2265 a_44916_1577# vss 0.0095f
C2266 a_47480_2002# vss 0.41829f
C2267 a_46620_1580# vss 0.52799f
C2268 a_47136_2122# vss 1.12757f
C2269 ShiftReg_row_10_2$1_0.DFF_2phase_1_2.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2270 a_42361_1539# vss 0.0072f
C2271 a_40748_1577# vss 0.0042f
C2272 a_41140_1577# vss 0.0095f
C2273 a_45016_2002# vss 0.42109f
C2274 a_44156_1580# vss 0.53063f
C2275 a_46152_1562# vss 1.18067f
C2276 a_44672_2122# vss 1.14287f
C2277 swmatrix_Tgate_0.gated_control vss 3.1994f
C2278 a_43688_1562# vss 1.1833f
C2279 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2280 ShiftReg_row_10_2$1_0.Q[7] vss 1.42957f
C2281 a_38284_1577# vss 0.0042f
C2282 a_38676_1577# vss 0.0095f
C2283 a_41240_2002# vss 0.41829f
C2284 a_40380_1580# vss 0.52799f
C2285 a_40896_2122# vss 1.12757f
C2286 ShiftReg_row_10_2$1_0.DFF_2phase_1_3.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2287 a_36121_1539# vss 0.0072f
C2288 a_34508_1577# vss 0.0042f
C2289 a_34900_1577# vss 0.0095f
C2290 a_38776_2002# vss 0.42109f
C2291 a_37916_1580# vss 0.53063f
C2292 a_39912_1562# vss 1.18067f
C2293 a_38432_2122# vss 1.14287f
C2294 swmatrix_Tgate_6.gated_control vss 3.1994f
C2295 a_37448_1562# vss 1.1833f
C2296 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2297 ShiftReg_row_10_2$1_0.Q[6] vss 1.42957f
C2298 a_32044_1577# vss 0.0042f
C2299 a_32436_1577# vss 0.0095f
C2300 a_35000_2002# vss 0.41829f
C2301 a_34140_1580# vss 0.52799f
C2302 a_34656_2122# vss 1.12757f
C2303 ShiftReg_row_10_2$1_0.DFF_2phase_1_4.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2304 a_29881_1539# vss 0.0072f
C2305 a_28268_1577# vss 0.0042f
C2306 a_28660_1577# vss 0.0095f
C2307 a_32536_2002# vss 0.42109f
C2308 a_31676_1580# vss 0.53063f
C2309 a_33672_1562# vss 1.18067f
C2310 a_32192_2122# vss 1.14287f
C2311 swmatrix_Tgate_5.gated_control vss 3.1994f
C2312 a_31208_1562# vss 1.1833f
C2313 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2314 ShiftReg_row_10_2$1_0.Q[5] vss 1.42957f
C2315 a_25804_1577# vss 0.0042f
C2316 a_26196_1577# vss 0.0095f
C2317 a_28760_2002# vss 0.41829f
C2318 a_27900_1580# vss 0.52799f
C2319 a_28416_2122# vss 1.12757f
C2320 ShiftReg_row_10_2$1_0.DFF_2phase_1_5.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2321 a_23641_1539# vss 0.0072f
C2322 a_22028_1577# vss 0.0042f
C2323 a_22420_1577# vss 0.0095f
C2324 a_26296_2002# vss 0.42109f
C2325 a_25436_1580# vss 0.53063f
C2326 a_27432_1562# vss 1.18067f
C2327 a_25952_2122# vss 1.14287f
C2328 swmatrix_Tgate_7.gated_control vss 3.1994f
C2329 a_24968_1562# vss 1.1833f
C2330 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2331 ShiftReg_row_10_2$1_0.Q[4] vss 1.42957f
C2332 a_19564_1577# vss 0.0042f
C2333 a_19956_1577# vss 0.0095f
C2334 a_22520_2002# vss 0.41829f
C2335 a_21660_1580# vss 0.52799f
C2336 a_22176_2122# vss 1.12757f
C2337 ShiftReg_row_10_2$1_0.DFF_2phase_1_6.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2338 a_17401_1539# vss 0.0072f
C2339 a_15788_1577# vss 0.0042f
C2340 a_16180_1577# vss 0.0095f
C2341 a_20056_2002# vss 0.42109f
C2342 a_19196_1580# vss 0.53063f
C2343 a_21192_1562# vss 1.18067f
C2344 a_19712_2122# vss 1.14287f
C2345 swmatrix_Tgate_4.gated_control vss 3.1994f
C2346 a_18728_1562# vss 1.1833f
C2347 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2348 ShiftReg_row_10_2$1_0.Q[3] vss 1.42957f
C2349 a_13324_1577# vss 0.0042f
C2350 a_13716_1577# vss 0.0095f
C2351 a_16280_2002# vss 0.41829f
C2352 a_15420_1580# vss 0.52799f
C2353 a_15936_2122# vss 1.12757f
C2354 ShiftReg_row_10_2$1_0.DFF_2phase_1_7.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2355 a_11161_1539# vss 0.0072f
C2356 a_9548_1577# vss 0.0042f
C2357 a_9940_1577# vss 0.0095f
C2358 a_13816_2002# vss 0.42109f
C2359 a_12956_1580# vss 0.53063f
C2360 a_14952_1562# vss 1.18067f
C2361 a_13472_2122# vss 1.14287f
C2362 swmatrix_Tgate_8.gated_control vss 3.20673f
C2363 a_12488_1562# vss 1.1833f
C2364 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.76917f
C2365 ShiftReg_row_10_2$1_0.Q[2] vss 1.42957f
C2366 a_7084_1577# vss 0.0042f
C2367 a_7476_1577# vss 0.0095f
C2368 a_10040_2002# vss 0.41829f
C2369 a_9180_1580# vss 0.52799f
C2370 a_9696_2122# vss 1.12757f
C2371 ShiftReg_row_10_2$1_0.DFF_2phase_1_9.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66671f
C2372 a_4921_1539# vss 0.0072f
C2373 a_3308_1577# vss 0.0042f
C2374 a_3700_1577# vss 0.0095f
C2375 a_7576_2002# vss 0.42109f
C2376 a_6716_1580# vss 0.53063f
C2377 a_8712_1562# vss 1.18067f
C2378 a_7232_2122# vss 1.14287f
C2379 swmatrix_Tgate_9.gated_control vss 3.24591f
C2380 a_6248_1562# vss 1.1833f
C2381 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__nand2_1_0.ZN vss 0.77126f
C2382 ShiftReg_row_10_2$1_0.Q[1] vss 1.43631f
C2383 a_844_1577# vss 0.0042f
C2384 a_1236_1577# vss 0.0095f
C2385 a_3800_2002# vss 0.4181f
C2386 a_2940_1580# vss 0.5278f
C2387 a_3456_2122# vss 1.12752f
C2388 ShiftReg_row_10_2$1_0.DFF_2phase_1_8.gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1.Q vss 0.66669f
C2389 a_1336_2002# vss 0.42132f
C2390 a_476_1580# vss 0.53083f
C2391 a_2472_1562# vss 1.18053f
C2392 a_992_2122# vss 1.1431f
C2393 a_8_1562# vss 1.19608f
C2394 BUS[10].t3 vss 0.08734f
C2395 BUS[10].t4 vss 0.08734f
C2396 BUS[10].n0 vss 0.4704f
C2397 BUS[10].t5 vss 0.08734f
C2398 BUS[10].t1 vss 0.08734f
C2399 BUS[10].n1 vss 0.46764f
C2400 BUS[10].n2 vss 0.27386f
C2401 BUS[10].t0 vss 0.08734f
C2402 BUS[10].t2 vss 0.08734f
C2403 BUS[10].n3 vss 0.46764f
C2404 BUS[10].n4 vss 0.23641f
C2405 BUS[10].t8 vss 0.08734f
C2406 BUS[10].t17 vss 0.08734f
C2407 BUS[10].n5 vss 0.47045f
C2408 BUS[10].n6 vss 0.20977f
C2409 BUS[10].t11 vss 0.08734f
C2410 BUS[10].t14 vss 0.08734f
C2411 BUS[10].n7 vss 0.47317f
C2412 BUS[10].t23 vss 0.08734f
C2413 BUS[10].t6 vss 0.08734f
C2414 BUS[10].n8 vss 0.47045f
C2415 BUS[10].n9 vss 0.26765f
C2416 BUS[10].t15 vss 0.08734f
C2417 BUS[10].t19 vss 0.08734f
C2418 BUS[10].n10 vss 0.47045f
C2419 BUS[10].n11 vss 0.15534f
C2420 BUS[10].t7 vss 0.08734f
C2421 BUS[10].t18 vss 0.08734f
C2422 BUS[10].n12 vss 0.47045f
C2423 BUS[10].n13 vss 0.15534f
C2424 BUS[10].t21 vss 0.08734f
C2425 BUS[10].t9 vss 0.08734f
C2426 BUS[10].n14 vss 0.47045f
C2427 BUS[10].n15 vss 0.15534f
C2428 BUS[10].t12 vss 0.08734f
C2429 BUS[10].t22 vss 0.08734f
C2430 BUS[10].n16 vss 0.47045f
C2431 BUS[10].n17 vss 0.15534f
C2432 BUS[10].t10 vss 0.08734f
C2433 BUS[10].t13 vss 0.08734f
C2434 BUS[10].n18 vss 0.47045f
C2435 BUS[10].n19 vss 0.15534f
C2436 BUS[10].t16 vss 0.08734f
C2437 BUS[10].t20 vss 0.08734f
C2438 BUS[10].n20 vss 0.47045f
C2439 BUS[10].n21 vss 0.10378f
C2440 BUS[10].n22 vss 0.3948f
C2441 BUS[3].t19 vss 0.08734f
C2442 BUS[3].t22 vss 0.08734f
C2443 BUS[3].n0 vss 0.4704f
C2444 BUS[3].t21 vss 0.08734f
C2445 BUS[3].t23 vss 0.08734f
C2446 BUS[3].n1 vss 0.46764f
C2447 BUS[3].n2 vss 0.27386f
C2448 BUS[3].t20 vss 0.08734f
C2449 BUS[3].t18 vss 0.08734f
C2450 BUS[3].n3 vss 0.46764f
C2451 BUS[3].n4 vss 0.23641f
C2452 BUS[3].t5 vss 0.08734f
C2453 BUS[3].t8 vss 0.08734f
C2454 BUS[3].n5 vss 0.47045f
C2455 BUS[3].n6 vss 0.20977f
C2456 BUS[3].t14 vss 0.08734f
C2457 BUS[3].t4 vss 0.08734f
C2458 BUS[3].n7 vss 0.47317f
C2459 BUS[3].t7 vss 0.08734f
C2460 BUS[3].t11 vss 0.08734f
C2461 BUS[3].n8 vss 0.47045f
C2462 BUS[3].n9 vss 0.26765f
C2463 BUS[3].t17 vss 0.08734f
C2464 BUS[3].t2 vss 0.08734f
C2465 BUS[3].n10 vss 0.47045f
C2466 BUS[3].n11 vss 0.15534f
C2467 BUS[3].t12 vss 0.08734f
C2468 BUS[3].t13 vss 0.08734f
C2469 BUS[3].n12 vss 0.47045f
C2470 BUS[3].n13 vss 0.15534f
C2471 BUS[3].t3 vss 0.08734f
C2472 BUS[3].t6 vss 0.08734f
C2473 BUS[3].n14 vss 0.47045f
C2474 BUS[3].n15 vss 0.15534f
C2475 BUS[3].t9 vss 0.08734f
C2476 BUS[3].t15 vss 0.08734f
C2477 BUS[3].n16 vss 0.47045f
C2478 BUS[3].n17 vss 0.15534f
C2479 BUS[3].t0 vss 0.08734f
C2480 BUS[3].t10 vss 0.08734f
C2481 BUS[3].n18 vss 0.47045f
C2482 BUS[3].n19 vss 0.15534f
C2483 BUS[3].t16 vss 0.08734f
C2484 BUS[3].t1 vss 0.08734f
C2485 BUS[3].n20 vss 0.47045f
C2486 BUS[3].n21 vss 0.10378f
C2487 BUS[3].n22 vss 0.3948f
C2488 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2489 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2490 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12308f
C2491 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2492 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2493 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C2494 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2495 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2496 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2497 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2498 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2499 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2500 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2501 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2502 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2503 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2504 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2505 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2506 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2507 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2508 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2509 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2510 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2511 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2512 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2513 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2514 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2515 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C2516 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2517 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C2518 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2519 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2520 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2521 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C2522 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2523 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2524 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2525 swmatrix_Tgate_4.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2526 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2527 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2528 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12308f
C2529 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2530 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2531 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2532 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2533 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C2534 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2535 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C2536 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2537 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C2538 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2539 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2540 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2541 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2542 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2543 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2544 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2545 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2546 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2547 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2548 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2549 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2550 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2551 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2552 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2553 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2554 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2555 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2556 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2557 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2558 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2559 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2560 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2561 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C2562 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2563 swmatrix_Tgate_8.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2564 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2565 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2566 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12308f
C2567 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2568 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2569 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2570 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2571 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2572 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2573 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2574 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2575 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2576 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2577 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2578 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2579 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2580 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2581 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2582 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2583 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2584 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2585 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2586 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2587 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C2588 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2589 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2590 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2591 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C2592 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2593 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C2594 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2595 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C2596 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2597 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2598 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2599 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2600 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2601 swmatrix_Tgate_2.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2602 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2603 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2604 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12308f
C2605 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2606 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2607 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2608 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2609 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2610 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2611 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C2612 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2613 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2614 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2615 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2616 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2617 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2618 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2619 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2620 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2621 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2622 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2623 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2624 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2625 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2626 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2627 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2628 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2629 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C2630 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2631 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2632 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2633 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C2634 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2635 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2636 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2637 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C2638 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2639 swmatrix_Tgate_1.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2640 PHI_1.t18 vss 0.12714f
C2641 PHI_1.t0 vss 0.0703f
C2642 PHI_1.n0 vss 0.1265f
C2643 PHI_1.t4 vss 0.12714f
C2644 PHI_1.t6 vss 0.0703f
C2645 PHI_1.n1 vss 0.1265f
C2646 PHI_1.n2 vss 1.47113f
C2647 PHI_1.t8 vss 0.12714f
C2648 PHI_1.t10 vss 0.0703f
C2649 PHI_1.n3 vss 0.1265f
C2650 PHI_1.n4 vss 1.47113f
C2651 PHI_1.t16 vss 0.12714f
C2652 PHI_1.t17 vss 0.0703f
C2653 PHI_1.n5 vss 0.1265f
C2654 PHI_1.n6 vss 1.47113f
C2655 PHI_1.t19 vss 0.12714f
C2656 PHI_1.t7 vss 0.0703f
C2657 PHI_1.n7 vss 0.1265f
C2658 PHI_1.n8 vss 1.47113f
C2659 PHI_1.t11 vss 0.12714f
C2660 PHI_1.t14 vss 0.0703f
C2661 PHI_1.n9 vss 0.1265f
C2662 PHI_1.n10 vss 1.47113f
C2663 PHI_1.t12 vss 0.12714f
C2664 PHI_1.t15 vss 0.0703f
C2665 PHI_1.n11 vss 0.1265f
C2666 PHI_1.n12 vss 1.47113f
C2667 PHI_1.t1 vss 0.12714f
C2668 PHI_1.t5 vss 0.0703f
C2669 PHI_1.n13 vss 0.1265f
C2670 PHI_1.n14 vss 1.47113f
C2671 PHI_1.t9 vss 0.12714f
C2672 PHI_1.t13 vss 0.0703f
C2673 PHI_1.n15 vss 0.1265f
C2674 PHI_1.n16 vss 1.47113f
C2675 PHI_1.t2 vss 0.12714f
C2676 PHI_1.t3 vss 0.0703f
C2677 PHI_1.n17 vss 0.1265f
C2678 PHI_1.n18 vss 1.47113f
C2679 enable.t1 vss 0.01609f
C2680 enable.t7 vss 0.01933f
C2681 enable.n0 vss 0.01817f
C2682 enable.n1 vss 0.00583f
C2683 enable.t13 vss 0.01609f
C2684 enable.t0 vss 0.01933f
C2685 enable.n2 vss 0.01817f
C2686 enable.n3 vss 0.00583f
C2687 enable.t9 vss 0.01609f
C2688 enable.t15 vss 0.01933f
C2689 enable.n4 vss 0.01817f
C2690 enable.n5 vss 0.00583f
C2691 enable.t16 vss 0.01609f
C2692 enable.t5 vss 0.01933f
C2693 enable.n6 vss 0.01817f
C2694 enable.n7 vss 0.00583f
C2695 enable.t12 vss 0.01609f
C2696 enable.t19 vss 0.01933f
C2697 enable.n8 vss 0.01817f
C2698 enable.n9 vss 0.00583f
C2699 enable.t6 vss 0.01609f
C2700 enable.t17 vss 0.01933f
C2701 enable.n10 vss 0.01817f
C2702 enable.n11 vss 0.00583f
C2703 enable.t18 vss 0.01609f
C2704 enable.t8 vss 0.01933f
C2705 enable.n12 vss 0.01817f
C2706 enable.n13 vss 0.00583f
C2707 enable.t14 vss 0.01609f
C2708 enable.t4 vss 0.01933f
C2709 enable.n14 vss 0.01817f
C2710 enable.n15 vss 0.00583f
C2711 enable.t3 vss 0.01609f
C2712 enable.t11 vss 0.01933f
C2713 enable.n16 vss 0.01817f
C2714 enable.n17 vss 0.00583f
C2715 enable.t2 vss 0.01609f
C2716 enable.t10 vss 0.01933f
C2717 enable.n18 vss 0.01817f
C2718 enable.n19 vss 0.11876f
C2719 enable.n20 vss 0.17899f
C2720 enable.n21 vss 0.17899f
C2721 enable.n22 vss 0.17899f
C2722 enable.n23 vss 0.17899f
C2723 enable.n24 vss 0.17899f
C2724 enable.n25 vss 0.17899f
C2725 enable.n26 vss 0.17899f
C2726 enable.n27 vss 0.17899f
C2727 enable.n28 vss 0.17899f
C2728 BUS[9].t9 vss 0.08734f
C2729 BUS[9].t10 vss 0.08734f
C2730 BUS[9].n0 vss 0.4704f
C2731 BUS[9].t12 vss 0.08734f
C2732 BUS[9].t14 vss 0.08734f
C2733 BUS[9].n1 vss 0.46764f
C2734 BUS[9].n2 vss 0.27386f
C2735 BUS[9].t13 vss 0.08734f
C2736 BUS[9].t11 vss 0.08734f
C2737 BUS[9].n3 vss 0.46764f
C2738 BUS[9].n4 vss 0.23641f
C2739 BUS[9].t15 vss 0.08734f
C2740 BUS[9].t5 vss 0.08734f
C2741 BUS[9].n5 vss 0.47045f
C2742 BUS[9].n6 vss 0.20977f
C2743 BUS[9].t18 vss 0.08734f
C2744 BUS[9].t0 vss 0.08734f
C2745 BUS[9].n7 vss 0.47317f
C2746 BUS[9].t1 vss 0.08734f
C2747 BUS[9].t21 vss 0.08734f
C2748 BUS[9].n8 vss 0.47045f
C2749 BUS[9].n9 vss 0.26765f
C2750 BUS[9].t8 vss 0.08734f
C2751 BUS[9].t23 vss 0.08734f
C2752 BUS[9].n10 vss 0.47045f
C2753 BUS[9].n11 vss 0.15534f
C2754 BUS[9].t3 vss 0.08734f
C2755 BUS[9].t4 vss 0.08734f
C2756 BUS[9].n12 vss 0.47045f
C2757 BUS[9].n13 vss 0.15534f
C2758 BUS[9].t16 vss 0.08734f
C2759 BUS[9].t2 vss 0.08734f
C2760 BUS[9].n14 vss 0.47045f
C2761 BUS[9].n15 vss 0.15534f
C2762 BUS[9].t19 vss 0.08734f
C2763 BUS[9].t20 vss 0.08734f
C2764 BUS[9].n16 vss 0.47045f
C2765 BUS[9].n17 vss 0.15534f
C2766 BUS[9].t7 vss 0.08734f
C2767 BUS[9].t22 vss 0.08734f
C2768 BUS[9].n18 vss 0.47045f
C2769 BUS[9].n19 vss 0.15534f
C2770 BUS[9].t6 vss 0.08734f
C2771 BUS[9].t17 vss 0.08734f
C2772 BUS[9].n20 vss 0.47045f
C2773 BUS[9].n21 vss 0.10378f
C2774 BUS[9].n22 vss 0.3948f
C2775 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2776 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2777 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12308f
C2778 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C2779 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2780 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2781 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2782 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2783 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2784 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2785 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2786 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2787 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2788 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C2789 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2790 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2791 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2792 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2793 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2794 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2795 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2796 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2797 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2798 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C2799 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2800 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2801 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2802 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2803 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2804 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2805 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2806 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2807 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2808 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2809 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2810 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C2811 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2812 swmatrix_Tgate_3.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2813 BUS[8].t5 vss 0.08734f
C2814 BUS[8].t9 vss 0.08734f
C2815 BUS[8].n0 vss 0.4704f
C2816 BUS[8].t8 vss 0.08734f
C2817 BUS[8].t10 vss 0.08734f
C2818 BUS[8].n1 vss 0.46764f
C2819 BUS[8].n2 vss 0.27386f
C2820 BUS[8].t6 vss 0.08734f
C2821 BUS[8].t7 vss 0.08734f
C2822 BUS[8].n3 vss 0.46764f
C2823 BUS[8].n4 vss 0.23641f
C2824 BUS[8].t12 vss 0.08734f
C2825 BUS[8].t14 vss 0.08734f
C2826 BUS[8].n5 vss 0.47045f
C2827 BUS[8].n6 vss 0.20977f
C2828 BUS[8].t20 vss 0.08734f
C2829 BUS[8].t1 vss 0.08734f
C2830 BUS[8].n7 vss 0.47317f
C2831 BUS[8].t0 vss 0.08734f
C2832 BUS[8].t23 vss 0.08734f
C2833 BUS[8].n8 vss 0.47045f
C2834 BUS[8].n9 vss 0.26765f
C2835 BUS[8].t19 vss 0.08734f
C2836 BUS[8].t16 vss 0.08734f
C2837 BUS[8].n10 vss 0.47045f
C2838 BUS[8].n11 vss 0.15534f
C2839 BUS[8].t11 vss 0.08734f
C2840 BUS[8].t2 vss 0.08734f
C2841 BUS[8].n12 vss 0.47045f
C2842 BUS[8].n13 vss 0.15534f
C2843 BUS[8].t15 vss 0.08734f
C2844 BUS[8].t3 vss 0.08734f
C2845 BUS[8].n14 vss 0.47045f
C2846 BUS[8].n15 vss 0.15534f
C2847 BUS[8].t21 vss 0.08734f
C2848 BUS[8].t22 vss 0.08734f
C2849 BUS[8].n16 vss 0.47045f
C2850 BUS[8].n17 vss 0.15534f
C2851 BUS[8].t18 vss 0.08734f
C2852 BUS[8].t13 vss 0.08734f
C2853 BUS[8].n18 vss 0.47045f
C2854 BUS[8].n19 vss 0.15534f
C2855 BUS[8].t4 vss 0.08734f
C2856 BUS[8].t17 vss 0.08734f
C2857 BUS[8].n20 vss 0.47045f
C2858 BUS[8].n21 vss 0.10378f
C2859 BUS[8].n22 vss 0.3948f
C2860 PHI_2.t18 vss 0.10988f
C2861 PHI_2.t1 vss 0.06075f
C2862 PHI_2.n0 vss 0.10937f
C2863 PHI_2.t4 vss 0.10988f
C2864 PHI_2.t11 vss 0.06075f
C2865 PHI_2.n1 vss 0.10937f
C2866 PHI_2.n2 vss 1.26325f
C2867 PHI_2.t15 vss 0.10988f
C2868 PHI_2.t17 vss 0.06075f
C2869 PHI_2.n3 vss 0.10937f
C2870 PHI_2.n4 vss 1.26325f
C2871 PHI_2.t0 vss 0.10988f
C2872 PHI_2.t3 vss 0.06075f
C2873 PHI_2.n5 vss 0.10937f
C2874 PHI_2.n6 vss 1.26325f
C2875 PHI_2.t6 vss 0.10988f
C2876 PHI_2.t7 vss 0.06075f
C2877 PHI_2.n7 vss 0.10937f
C2878 PHI_2.n8 vss 1.26325f
C2879 PHI_2.t12 vss 0.10988f
C2880 PHI_2.t14 vss 0.06075f
C2881 PHI_2.n9 vss 0.10937f
C2882 PHI_2.n10 vss 1.26325f
C2883 PHI_2.t16 vss 0.10988f
C2884 PHI_2.t5 vss 0.06075f
C2885 PHI_2.n11 vss 0.10937f
C2886 PHI_2.n12 vss 1.26325f
C2887 PHI_2.t8 vss 0.10988f
C2888 PHI_2.t10 vss 0.06075f
C2889 PHI_2.n13 vss 0.10937f
C2890 PHI_2.n14 vss 1.26325f
C2891 PHI_2.t9 vss 0.10988f
C2892 PHI_2.t13 vss 0.06075f
C2893 PHI_2.n15 vss 0.10937f
C2894 PHI_2.n16 vss 1.26325f
C2895 PHI_2.t19 vss 0.10988f
C2896 PHI_2.t2 vss 0.06075f
C2897 PHI_2.n17 vss 0.10937f
C2898 PHI_2.n18 vss 1.26325f
C2899 BUS[4].t19 vss 0.08734f
C2900 BUS[4].t21 vss 0.08734f
C2901 BUS[4].n0 vss 0.4704f
C2902 BUS[4].t20 vss 0.08734f
C2903 BUS[4].t23 vss 0.08734f
C2904 BUS[4].n1 vss 0.46764f
C2905 BUS[4].n2 vss 0.27386f
C2906 BUS[4].t22 vss 0.08734f
C2907 BUS[4].t18 vss 0.08734f
C2908 BUS[4].n3 vss 0.46764f
C2909 BUS[4].n4 vss 0.23641f
C2910 BUS[4].t15 vss 0.08734f
C2911 BUS[4].t1 vss 0.08734f
C2912 BUS[4].n5 vss 0.47045f
C2913 BUS[4].n6 vss 0.20977f
C2914 BUS[4].t7 vss 0.08734f
C2915 BUS[4].t9 vss 0.08734f
C2916 BUS[4].n7 vss 0.47317f
C2917 BUS[4].t0 vss 0.08734f
C2918 BUS[4].t8 vss 0.08734f
C2919 BUS[4].n8 vss 0.47045f
C2920 BUS[4].n9 vss 0.26765f
C2921 BUS[4].t10 vss 0.08734f
C2922 BUS[4].t13 vss 0.08734f
C2923 BUS[4].n10 vss 0.47045f
C2924 BUS[4].n11 vss 0.15534f
C2925 BUS[4].t16 vss 0.08734f
C2926 BUS[4].t5 vss 0.08734f
C2927 BUS[4].n12 vss 0.47045f
C2928 BUS[4].n13 vss 0.15534f
C2929 BUS[4].t14 vss 0.08734f
C2930 BUS[4].t17 vss 0.08734f
C2931 BUS[4].n14 vss 0.47045f
C2932 BUS[4].n15 vss 0.15534f
C2933 BUS[4].t6 vss 0.08734f
C2934 BUS[4].t3 vss 0.08734f
C2935 BUS[4].n16 vss 0.47045f
C2936 BUS[4].n17 vss 0.15534f
C2937 BUS[4].t11 vss 0.08734f
C2938 BUS[4].t2 vss 0.08734f
C2939 BUS[4].n18 vss 0.47045f
C2940 BUS[4].n19 vss 0.15534f
C2941 BUS[4].t4 vss 0.08734f
C2942 BUS[4].t12 vss 0.08734f
C2943 BUS[4].n20 vss 0.47045f
C2944 BUS[4].n21 vss 0.10378f
C2945 BUS[4].n22 vss 0.3948f
C2946 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C2947 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C2948 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12308f
C2949 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C2950 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C2951 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C2952 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C2953 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C2954 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C2955 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C2956 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C2957 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C2958 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C2959 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C2960 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C2961 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C2962 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C2963 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C2964 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C2965 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C2966 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C2967 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C2968 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C2969 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C2970 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C2971 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C2972 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C2973 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C2974 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C2975 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C2976 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C2977 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C2978 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C2979 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C2980 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C2981 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C2982 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C2983 swmatrix_Tgate_7.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C2984 BUS[6].t5 vss 0.08734f
C2985 BUS[6].t0 vss 0.08734f
C2986 BUS[6].n0 vss 0.4704f
C2987 BUS[6].t1 vss 0.08734f
C2988 BUS[6].t3 vss 0.08734f
C2989 BUS[6].n1 vss 0.46764f
C2990 BUS[6].n2 vss 0.27386f
C2991 BUS[6].t2 vss 0.08734f
C2992 BUS[6].t4 vss 0.08734f
C2993 BUS[6].n3 vss 0.46764f
C2994 BUS[6].n4 vss 0.23641f
C2995 BUS[6].t19 vss 0.08734f
C2996 BUS[6].t21 vss 0.08734f
C2997 BUS[6].n5 vss 0.47045f
C2998 BUS[6].n6 vss 0.20977f
C2999 BUS[6].t10 vss 0.08734f
C3000 BUS[6].t14 vss 0.08734f
C3001 BUS[6].n7 vss 0.47317f
C3002 BUS[6].t17 vss 0.08734f
C3003 BUS[6].t6 vss 0.08734f
C3004 BUS[6].n8 vss 0.47045f
C3005 BUS[6].n9 vss 0.26765f
C3006 BUS[6].t8 vss 0.08734f
C3007 BUS[6].t18 vss 0.08734f
C3008 BUS[6].n10 vss 0.47045f
C3009 BUS[6].n11 vss 0.15534f
C3010 BUS[6].t7 vss 0.08734f
C3011 BUS[6].t9 vss 0.08734f
C3012 BUS[6].n12 vss 0.47045f
C3013 BUS[6].n13 vss 0.15534f
C3014 BUS[6].t12 vss 0.08734f
C3015 BUS[6].t15 vss 0.08734f
C3016 BUS[6].n14 vss 0.47045f
C3017 BUS[6].n15 vss 0.15534f
C3018 BUS[6].t22 vss 0.08734f
C3019 BUS[6].t13 vss 0.08734f
C3020 BUS[6].n16 vss 0.47045f
C3021 BUS[6].n17 vss 0.15534f
C3022 BUS[6].t16 vss 0.08734f
C3023 BUS[6].t23 vss 0.08734f
C3024 BUS[6].n18 vss 0.47045f
C3025 BUS[6].n19 vss 0.15534f
C3026 BUS[6].t20 vss 0.08734f
C3027 BUS[6].t11 vss 0.08734f
C3028 BUS[6].n20 vss 0.47045f
C3029 BUS[6].n21 vss 0.10378f
C3030 BUS[6].n22 vss 0.3948f
C3031 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C3032 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C3033 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12308f
C3034 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C3035 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C3036 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C3037 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C3038 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C3039 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C3040 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C3041 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C3042 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C3043 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C3044 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C3045 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C3046 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C3047 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C3048 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C3049 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C3050 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C3051 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C3052 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C3053 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C3054 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C3055 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C3056 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C3057 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C3058 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C3059 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C3060 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C3061 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C3062 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C3063 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C3064 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C3065 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C3066 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C3067 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C3068 swmatrix_Tgate_6.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C3069 BUS[5].t3 vss 0.08734f
C3070 BUS[5].t1 vss 0.08734f
C3071 BUS[5].n0 vss 0.4704f
C3072 BUS[5].t2 vss 0.08734f
C3073 BUS[5].t5 vss 0.08734f
C3074 BUS[5].n1 vss 0.46764f
C3075 BUS[5].n2 vss 0.27386f
C3076 BUS[5].t4 vss 0.08734f
C3077 BUS[5].t0 vss 0.08734f
C3078 BUS[5].n3 vss 0.46764f
C3079 BUS[5].n4 vss 0.23641f
C3080 BUS[5].t6 vss 0.08734f
C3081 BUS[5].t14 vss 0.08734f
C3082 BUS[5].n5 vss 0.47045f
C3083 BUS[5].n6 vss 0.20977f
C3084 BUS[5].t11 vss 0.08734f
C3085 BUS[5].t19 vss 0.08734f
C3086 BUS[5].n7 vss 0.47317f
C3087 BUS[5].t9 vss 0.08734f
C3088 BUS[5].t12 vss 0.08734f
C3089 BUS[5].n8 vss 0.47045f
C3090 BUS[5].n9 vss 0.26765f
C3091 BUS[5].t20 vss 0.08734f
C3092 BUS[5].t22 vss 0.08734f
C3093 BUS[5].n10 vss 0.47045f
C3094 BUS[5].n11 vss 0.15534f
C3095 BUS[5].t7 vss 0.08734f
C3096 BUS[5].t15 vss 0.08734f
C3097 BUS[5].n12 vss 0.47045f
C3098 BUS[5].n13 vss 0.15534f
C3099 BUS[5].t17 vss 0.08734f
C3100 BUS[5].t8 vss 0.08734f
C3101 BUS[5].n14 vss 0.47045f
C3102 BUS[5].n15 vss 0.15534f
C3103 BUS[5].t10 vss 0.08734f
C3104 BUS[5].t18 vss 0.08734f
C3105 BUS[5].n16 vss 0.47045f
C3106 BUS[5].n17 vss 0.15534f
C3107 BUS[5].t21 vss 0.08734f
C3108 BUS[5].t23 vss 0.08734f
C3109 BUS[5].n18 vss 0.47045f
C3110 BUS[5].n19 vss 0.15534f
C3111 BUS[5].t13 vss 0.08734f
C3112 BUS[5].t16 vss 0.08734f
C3113 BUS[5].n20 vss 0.47045f
C3114 BUS[5].n21 vss 0.10378f
C3115 BUS[5].n22 vss 0.3948f
C3116 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C3117 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C3118 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12308f
C3119 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C3120 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C3121 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C3122 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C3123 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C3124 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C3125 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C3126 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C3127 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C3128 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C3129 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C3130 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C3131 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C3132 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C3133 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C3134 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C3135 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C3136 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C3137 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C3138 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C3139 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C3140 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C3141 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C3142 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C3143 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C3144 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C3145 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C3146 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C3147 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C3148 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C3149 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C3150 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C3151 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C3152 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C3153 swmatrix_Tgate_5.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C3154 BUS[1].t19 vss 0.08731f
C3155 BUS[1].t20 vss 0.08731f
C3156 BUS[1].n0 vss 0.47019f
C3157 BUS[1].t21 vss 0.08731f
C3158 BUS[1].t23 vss 0.08731f
C3159 BUS[1].n1 vss 0.46743f
C3160 BUS[1].n2 vss 0.27374f
C3161 BUS[1].t22 vss 0.08731f
C3162 BUS[1].t18 vss 0.08731f
C3163 BUS[1].n3 vss 0.46743f
C3164 BUS[1].n4 vss 0.2363f
C3165 BUS[1].t0 vss 0.08731f
C3166 BUS[1].t3 vss 0.08731f
C3167 BUS[1].n5 vss 0.47023f
C3168 BUS[1].n6 vss 0.20967f
C3169 BUS[1].t6 vss 0.08731f
C3170 BUS[1].t13 vss 0.08731f
C3171 BUS[1].n7 vss 0.47295f
C3172 BUS[1].t15 vss 0.08731f
C3173 BUS[1].t7 vss 0.08731f
C3174 BUS[1].n8 vss 0.47023f
C3175 BUS[1].n9 vss 0.26753f
C3176 BUS[1].t8 vss 0.08731f
C3177 BUS[1].t16 vss 0.08731f
C3178 BUS[1].n10 vss 0.47023f
C3179 BUS[1].n11 vss 0.15527f
C3180 BUS[1].t1 vss 0.08731f
C3181 BUS[1].t4 vss 0.08731f
C3182 BUS[1].n12 vss 0.47023f
C3183 BUS[1].n13 vss 0.15527f
C3184 BUS[1].t11 vss 0.08731f
C3185 BUS[1].t14 vss 0.08731f
C3186 BUS[1].n14 vss 0.47023f
C3187 BUS[1].n15 vss 0.15527f
C3188 BUS[1].t5 vss 0.08731f
C3189 BUS[1].t12 vss 0.08731f
C3190 BUS[1].n16 vss 0.47023f
C3191 BUS[1].n17 vss 0.15527f
C3192 BUS[1].t9 vss 0.08731f
C3193 BUS[1].t17 vss 0.08731f
C3194 BUS[1].n18 vss 0.47023f
C3195 BUS[1].n19 vss 0.15527f
C3196 BUS[1].t2 vss 0.08731f
C3197 BUS[1].t10 vss 0.08731f
C3198 BUS[1].n20 vss 0.47023f
C3199 BUS[1].n21 vss 0.10373f
C3200 BUS[1].n22 vss 0.39702f
C3201 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.06869f
C3202 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.09485f
C3203 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12308f
C3204 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C3205 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C3206 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C3207 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C3208 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C3209 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C3210 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C3211 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C3212 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C3213 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C3214 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C3215 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C3216 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C3217 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C3218 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C3219 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C3220 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C3221 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C3222 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C3223 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C3224 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C3225 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C3226 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C3227 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C3228 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12285f
C3229 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C3230 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C3231 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C3232 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C3233 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C3234 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C3235 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C3236 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C3237 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C3238 swmatrix_Tgate_9.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
C3239 BUS[2].t17 vss 0.08734f
C3240 BUS[2].t20 vss 0.08734f
C3241 BUS[2].n0 vss 0.4704f
C3242 BUS[2].t19 vss 0.08734f
C3243 BUS[2].t16 vss 0.08734f
C3244 BUS[2].n1 vss 0.46764f
C3245 BUS[2].n2 vss 0.27386f
C3246 BUS[2].t21 vss 0.08734f
C3247 BUS[2].t18 vss 0.08734f
C3248 BUS[2].n3 vss 0.46764f
C3249 BUS[2].n4 vss 0.23641f
C3250 BUS[2].t4 vss 0.08734f
C3251 BUS[2].t11 vss 0.08734f
C3252 BUS[2].n5 vss 0.47045f
C3253 BUS[2].n6 vss 0.20977f
C3254 BUS[2].t22 vss 0.08734f
C3255 BUS[2].t5 vss 0.08734f
C3256 BUS[2].n7 vss 0.47317f
C3257 BUS[2].t12 vss 0.08734f
C3258 BUS[2].t9 vss 0.08734f
C3259 BUS[2].n8 vss 0.47045f
C3260 BUS[2].n9 vss 0.26765f
C3261 BUS[2].t14 vss 0.08734f
C3262 BUS[2].t7 vss 0.08734f
C3263 BUS[2].n10 vss 0.47045f
C3264 BUS[2].n11 vss 0.15534f
C3265 BUS[2].t3 vss 0.08734f
C3266 BUS[2].t23 vss 0.08734f
C3267 BUS[2].n12 vss 0.47045f
C3268 BUS[2].n13 vss 0.15534f
C3269 BUS[2].t0 vss 0.08734f
C3270 BUS[2].t1 vss 0.08734f
C3271 BUS[2].n14 vss 0.47045f
C3272 BUS[2].n15 vss 0.15534f
C3273 BUS[2].t10 vss 0.08734f
C3274 BUS[2].t15 vss 0.08734f
C3275 BUS[2].n16 vss 0.47045f
C3276 BUS[2].n17 vss 0.15534f
C3277 BUS[2].t13 vss 0.08734f
C3278 BUS[2].t6 vss 0.08734f
C3279 BUS[2].n18 vss 0.47045f
C3280 BUS[2].n19 vss 0.15534f
C3281 BUS[2].t2 vss 0.08734f
C3282 BUS[2].t8 vss 0.08734f
C3283 BUS[2].n20 vss 0.47045f
C3284 BUS[2].n21 vss 0.10378f
C3285 BUS[2].n22 vss 0.3948f
C3286 vdd.t54 vss 0.00786f
C3287 vdd.t288 vss 0.00385f
C3288 vdd.n0 vss 0.0167f
C3289 vdd.t294 vss 0.0098f
C3290 vdd.t117 vss 0.00522f
C3291 vdd.t5 vss 0.00522f
C3292 vdd.n1 vss 0.01114f
C3293 vdd.t115 vss 0.0198f
C3294 vdd.t287 vss 0.08979f
C3295 vdd.t53 vss 0.14646f
C3296 vdd.t293 vss 0.12034f
C3297 vdd.t52 vss 0.08209f
C3298 vdd.t23 vss 0.10355f
C3299 vdd.t4 vss 0.10355f
C3300 vdd.t116 vss 0.14739f
C3301 vdd.t114 vss 0.17025f
C3302 vdd.n2 vss 0.10679f
C3303 vdd.t113 vss 0.00786f
C3304 vdd.t524 vss 0.00385f
C3305 vdd.n3 vss 0.0167f
C3306 vdd.t156 vss 0.0098f
C3307 vdd.t184 vss 0.00522f
C3308 vdd.t7 vss 0.00522f
C3309 vdd.n4 vss 0.01114f
C3310 vdd.t186 vss 0.0198f
C3311 vdd.t89 vss 0.01707f
C3312 vdd.t509 vss 0.01684f
C3313 vdd.t470 vss 0.01948f
C3314 vdd.t523 vss 0.08979f
C3315 vdd.t112 vss 0.14646f
C3316 vdd.t155 vss 0.12034f
C3317 vdd.t111 vss 0.08209f
C3318 vdd.t134 vss 0.10355f
C3319 vdd.t6 vss 0.10355f
C3320 vdd.t183 vss 0.14739f
C3321 vdd.t185 vss 0.16115f
C3322 vdd.t88 vss 0.0723f
C3323 vdd.t508 vss 0.10588f
C3324 vdd.t469 vss 0.11358f
C3325 vdd.n5 vss 0.14854f
C3326 vdd.n6 vss 0.10726f
C3327 vdd.t41 vss 0.00786f
C3328 vdd.t284 vss 0.00385f
C3329 vdd.n7 vss 0.0167f
C3330 vdd.t87 vss 0.0098f
C3331 vdd.t443 vss 0.00522f
C3332 vdd.t429 vss 0.00522f
C3333 vdd.n8 vss 0.01114f
C3334 vdd.t441 vss 0.0198f
C3335 vdd.t283 vss 0.08979f
C3336 vdd.t40 vss 0.14646f
C3337 vdd.t86 vss 0.12034f
C3338 vdd.t42 vss 0.08209f
C3339 vdd.t454 vss 0.10355f
C3340 vdd.t428 vss 0.10355f
C3341 vdd.t442 vss 0.14739f
C3342 vdd.t440 vss 0.17025f
C3343 vdd.n9 vss 0.10679f
C3344 vdd.t383 vss 0.00786f
C3345 vdd.t257 vss 0.00385f
C3346 vdd.n10 vss 0.0167f
C3347 vdd.t150 vss 0.0098f
C3348 vdd.t93 vss 0.00522f
C3349 vdd.t152 vss 0.00522f
C3350 vdd.n11 vss 0.01114f
C3351 vdd.t95 vss 0.0198f
C3352 vdd.t447 vss 0.01707f
C3353 vdd.t234 vss 0.01684f
C3354 vdd.t243 vss 0.01948f
C3355 vdd.t256 vss 0.08979f
C3356 vdd.t382 vss 0.14646f
C3357 vdd.t149 vss 0.12034f
C3358 vdd.t381 vss 0.08209f
C3359 vdd.t148 vss 0.10355f
C3360 vdd.t151 vss 0.10355f
C3361 vdd.t92 vss 0.14739f
C3362 vdd.t94 vss 0.16115f
C3363 vdd.t446 vss 0.0723f
C3364 vdd.t233 vss 0.10588f
C3365 vdd.t242 vss 0.11358f
C3366 vdd.n12 vss 0.14854f
C3367 vdd.n13 vss 0.10726f
C3368 vdd.t66 vss 0.00786f
C3369 vdd.t286 vss 0.00385f
C3370 vdd.n14 vss 0.0167f
C3371 vdd.t445 vss 0.0098f
C3372 vdd.t410 vss 0.00522f
C3373 vdd.t59 vss 0.00522f
C3374 vdd.n15 vss 0.01114f
C3375 vdd.t412 vss 0.0198f
C3376 vdd.t285 vss 0.08979f
C3377 vdd.t65 vss 0.14646f
C3378 vdd.t444 vss 0.12034f
C3379 vdd.t67 vss 0.08209f
C3380 vdd.t191 vss 0.10355f
C3381 vdd.t58 vss 0.10355f
C3382 vdd.t409 vss 0.14739f
C3383 vdd.t411 vss 0.17025f
C3384 vdd.n16 vss 0.10679f
C3385 vdd.t271 vss 0.00786f
C3386 vdd.t255 vss 0.00385f
C3387 vdd.n17 vss 0.0167f
C3388 vdd.t371 vss 0.0098f
C3389 vdd.t435 vss 0.00522f
C3390 vdd.t373 vss 0.00522f
C3391 vdd.n18 vss 0.01114f
C3392 vdd.t437 vss 0.0198f
C3393 vdd.t165 vss 0.01707f
C3394 vdd.t190 vss 0.01684f
C3395 vdd.t97 vss 0.01948f
C3396 vdd.t254 vss 0.08979f
C3397 vdd.t270 vss 0.14646f
C3398 vdd.t370 vss 0.12034f
C3399 vdd.t269 vss 0.08209f
C3400 vdd.t125 vss 0.10355f
C3401 vdd.t372 vss 0.10355f
C3402 vdd.t434 vss 0.14739f
C3403 vdd.t436 vss 0.16115f
C3404 vdd.t164 vss 0.0723f
C3405 vdd.t189 vss 0.10588f
C3406 vdd.t96 vss 0.11358f
C3407 vdd.n19 vss 0.14854f
C3408 vdd.n20 vss 0.10726f
C3409 vdd.t161 vss 0.00786f
C3410 vdd.t307 vss 0.00385f
C3411 vdd.n21 vss 0.0167f
C3412 vdd.t167 vss 0.0098f
C3413 vdd.t536 vss 0.00522f
C3414 vdd.t182 vss 0.00522f
C3415 vdd.n22 vss 0.01114f
C3416 vdd.t534 vss 0.0198f
C3417 vdd.t306 vss 0.08979f
C3418 vdd.t160 vss 0.14646f
C3419 vdd.t166 vss 0.12034f
C3420 vdd.t159 vss 0.08209f
C3421 vdd.t387 vss 0.10355f
C3422 vdd.t181 vss 0.10355f
C3423 vdd.t535 vss 0.14739f
C3424 vdd.t533 vss 0.17025f
C3425 vdd.n23 vss 0.10679f
C3426 vdd.t30 vss 0.00786f
C3427 vdd.t520 vss 0.00385f
C3428 vdd.n24 vss 0.0167f
C3429 vdd.t170 vss 0.0098f
C3430 vdd.t460 vss 0.00522f
C3431 vdd.t120 vss 0.00522f
C3432 vdd.n25 vss 0.01114f
C3433 vdd.t462 vss 0.0198f
C3434 vdd.t407 vss 0.01707f
C3435 vdd.t1 vss 0.01684f
C3436 vdd.t37 vss 0.01948f
C3437 vdd.t519 vss 0.08979f
C3438 vdd.t29 vss 0.14646f
C3439 vdd.t169 vss 0.12034f
C3440 vdd.t28 vss 0.08209f
C3441 vdd.t374 vss 0.10355f
C3442 vdd.t119 vss 0.10355f
C3443 vdd.t459 vss 0.14739f
C3444 vdd.t461 vss 0.16115f
C3445 vdd.t406 vss 0.0723f
C3446 vdd.t0 vss 0.10588f
C3447 vdd.t36 vss 0.11358f
C3448 vdd.n26 vss 0.14854f
C3449 vdd.n27 vss 0.10726f
C3450 vdd.t515 vss 0.00786f
C3451 vdd.t305 vss 0.00385f
C3452 vdd.n28 vss 0.0167f
C3453 vdd.t405 vss 0.0098f
C3454 vdd.t456 vss 0.00522f
C3455 vdd.t476 vss 0.00522f
C3456 vdd.n29 vss 0.01114f
C3457 vdd.t458 vss 0.0198f
C3458 vdd.t304 vss 0.08979f
C3459 vdd.t514 vss 0.14646f
C3460 vdd.t404 vss 0.12034f
C3461 vdd.t516 vss 0.08209f
C3462 vdd.t147 vss 0.10355f
C3463 vdd.t475 vss 0.10355f
C3464 vdd.t455 vss 0.14739f
C3465 vdd.t457 vss 0.17025f
C3466 vdd.n30 vss 0.10679f
C3467 vdd.t482 vss 0.00786f
C3468 vdd.t526 vss 0.00385f
C3469 vdd.n31 vss 0.0167f
C3470 vdd.t127 vss 0.0098f
C3471 vdd.t424 vss 0.00522f
C3472 vdd.t99 vss 0.00522f
C3473 vdd.n32 vss 0.01114f
C3474 vdd.t426 vss 0.0198f
C3475 vdd.t133 vss 0.01707f
C3476 vdd.t232 vss 0.01684f
C3477 vdd.t12 vss 0.01948f
C3478 vdd.t525 vss 0.08979f
C3479 vdd.t481 vss 0.14646f
C3480 vdd.t126 vss 0.12034f
C3481 vdd.t483 vss 0.08209f
C3482 vdd.t168 vss 0.10355f
C3483 vdd.t98 vss 0.10355f
C3484 vdd.t423 vss 0.14739f
C3485 vdd.t425 vss 0.16115f
C3486 vdd.t132 vss 0.0723f
C3487 vdd.t231 vss 0.10588f
C3488 vdd.t11 vss 0.11358f
C3489 vdd.n33 vss 0.14854f
C3490 vdd.n34 vss 0.10726f
C3491 vdd.t141 vss 0.00786f
C3492 vdd.t336 vss 0.00385f
C3493 vdd.n35 vss 0.0167f
C3494 vdd.t131 vss 0.0098f
C3495 vdd.t318 vss 0.00522f
C3496 vdd.t176 vss 0.00522f
C3497 vdd.n36 vss 0.01114f
C3498 vdd.t320 vss 0.0198f
C3499 vdd.t335 vss 0.08979f
C3500 vdd.t140 vss 0.14646f
C3501 vdd.t130 vss 0.12034f
C3502 vdd.t142 vss 0.08209f
C3503 vdd.t100 vss 0.10355f
C3504 vdd.t175 vss 0.10355f
C3505 vdd.t317 vss 0.14739f
C3506 vdd.t319 vss 0.17025f
C3507 vdd.n37 vss 0.10679f
C3508 vdd.t323 vss 0.00786f
C3509 vdd.t34 vss 0.00385f
C3510 vdd.n38 vss 0.0167f
C3511 vdd.t340 vss 0.0098f
C3512 vdd.t144 vss 0.00522f
C3513 vdd.t449 vss 0.00522f
C3514 vdd.n39 vss 0.01114f
C3515 vdd.t146 vss 0.0198f
C3516 vdd.t178 vss 0.01707f
C3517 vdd.t39 vss 0.01684f
C3518 vdd.t51 vss 0.01948f
C3519 vdd.t33 vss 0.08979f
C3520 vdd.t322 vss 0.14646f
C3521 vdd.t339 vss 0.12034f
C3522 vdd.t321 vss 0.08209f
C3523 vdd.t153 vss 0.10355f
C3524 vdd.t448 vss 0.10355f
C3525 vdd.t143 vss 0.14739f
C3526 vdd.t145 vss 0.16115f
C3527 vdd.t177 vss 0.0723f
C3528 vdd.t38 vss 0.10588f
C3529 vdd.t50 vss 0.11358f
C3530 vdd.n40 vss 0.14854f
C3531 vdd.n41 vss 0.10726f
C3532 vdd.t265 vss 0.00786f
C3533 vdd.t273 vss 0.00385f
C3534 vdd.n42 vss 0.0167f
C3535 vdd.t180 vss 0.0098f
C3536 vdd.t366 vss 0.00522f
C3537 vdd.t414 vss 0.00522f
C3538 vdd.n43 vss 0.01114f
C3539 vdd.t364 vss 0.0198f
C3540 vdd.t272 vss 0.08979f
C3541 vdd.t264 vss 0.14646f
C3542 vdd.t179 vss 0.12034f
C3543 vdd.t266 vss 0.08209f
C3544 vdd.t316 vss 0.10355f
C3545 vdd.t413 vss 0.10355f
C3546 vdd.t365 vss 0.14739f
C3547 vdd.t363 vss 0.17025f
C3548 vdd.n44 vss 0.10679f
C3549 vdd.t369 vss 0.00786f
C3550 vdd.t224 vss 0.00385f
C3551 vdd.n45 vss 0.0167f
C3552 vdd.t110 vss 0.0098f
C3553 vdd.t495 vss 0.00522f
C3554 vdd.t158 vss 0.00522f
C3555 vdd.n46 vss 0.01114f
C3556 vdd.t493 vss 0.0198f
C3557 vdd.t453 vss 0.01707f
C3558 vdd.t3 vss 0.01684f
C3559 vdd.t268 vss 0.01948f
C3560 vdd.t223 vss 0.08979f
C3561 vdd.t368 vss 0.14646f
C3562 vdd.t109 vss 0.12034f
C3563 vdd.t367 vss 0.08209f
C3564 vdd.t35 vss 0.10355f
C3565 vdd.t157 vss 0.10355f
C3566 vdd.t494 vss 0.14739f
C3567 vdd.t492 vss 0.16115f
C3568 vdd.t452 vss 0.0723f
C3569 vdd.t2 vss 0.10588f
C3570 vdd.t267 vss 0.11358f
C3571 vdd.n47 vss 0.14854f
C3572 vdd.n48 vss 0.10726f
C3573 vdd.t193 vss 0.00786f
C3574 vdd.t282 vss 0.00385f
C3575 vdd.n49 vss 0.0167f
C3576 vdd.t451 vss 0.0098f
C3577 vdd.t16 vss 0.00522f
C3578 vdd.t380 vss 0.00522f
C3579 vdd.n50 vss 0.01114f
C3580 vdd.t14 vss 0.0198f
C3581 vdd.t281 vss 0.08979f
C3582 vdd.t192 vss 0.14646f
C3583 vdd.t450 vss 0.12034f
C3584 vdd.t194 vss 0.08209f
C3585 vdd.t44 vss 0.10355f
C3586 vdd.t379 vss 0.10355f
C3587 vdd.t15 vss 0.14739f
C3588 vdd.t13 vss 0.17025f
C3589 vdd.n51 vss 0.10679f
C3590 vdd.t48 vss 0.00786f
C3591 vdd.t528 vss 0.00385f
C3592 vdd.n52 vss 0.0167f
C3593 vdd.t27 vss 0.0098f
C3594 vdd.t124 vss 0.00522f
C3595 vdd.t490 vss 0.00522f
C3596 vdd.n53 vss 0.01114f
C3597 vdd.t122 vss 0.0198f
C3598 vdd.t174 vss 0.01707f
C3599 vdd.t56 vss 0.01684f
C3600 vdd.t91 vss 0.01948f
C3601 vdd.t527 vss 0.08979f
C3602 vdd.t47 vss 0.14646f
C3603 vdd.t26 vss 0.12034f
C3604 vdd.t49 vss 0.08209f
C3605 vdd.t139 vss 0.10355f
C3606 vdd.t489 vss 0.10355f
C3607 vdd.t123 vss 0.14739f
C3608 vdd.t121 vss 0.16115f
C3609 vdd.t173 vss 0.0723f
C3610 vdd.t55 vss 0.10588f
C3611 vdd.t90 vss 0.11358f
C3612 vdd.n54 vss 0.14854f
C3613 vdd.n55 vss 0.10726f
C3614 vdd.t386 vss 0.00786f
C3615 vdd.t280 vss 0.00385f
C3616 vdd.n56 vss 0.0167f
C3617 vdd.t172 vss 0.0098f
C3618 vdd.t102 vss 0.00522f
C3619 vdd.t518 vss 0.00522f
C3620 vdd.n57 vss 0.01114f
C3621 vdd.t104 vss 0.0198f
C3622 vdd.t279 vss 0.08979f
C3623 vdd.t385 vss 0.14646f
C3624 vdd.t171 vss 0.12034f
C3625 vdd.t384 vss 0.08209f
C3626 vdd.t427 vss 0.10355f
C3627 vdd.t517 vss 0.10355f
C3628 vdd.t101 vss 0.14739f
C3629 vdd.t103 vss 0.17025f
C3630 vdd.n58 vss 0.10679f
C3631 vdd.t196 vss 0.00786f
C3632 vdd.t32 vss 0.00385f
C3633 vdd.n59 vss 0.0167f
C3634 vdd.t106 vss 0.0098f
C3635 vdd.t472 vss 0.00522f
C3636 vdd.t263 vss 0.00522f
C3637 vdd.n60 vss 0.01114f
C3638 vdd.t474 vss 0.0198f
C3639 vdd.t419 vss 0.01707f
C3640 vdd.t513 vss 0.01684f
C3641 vdd.t290 vss 0.01948f
C3642 vdd.t31 vss 0.08979f
C3643 vdd.t195 vss 0.14646f
C3644 vdd.t105 vss 0.12034f
C3645 vdd.t197 vss 0.08209f
C3646 vdd.t315 vss 0.10355f
C3647 vdd.t262 vss 0.10355f
C3648 vdd.t471 vss 0.14739f
C3649 vdd.t473 vss 0.16115f
C3650 vdd.t418 vss 0.0723f
C3651 vdd.t512 vss 0.10588f
C3652 vdd.t289 vss 0.11358f
C3653 vdd.n61 vss 0.14854f
C3654 vdd.n62 vss 0.10726f
C3655 vdd.t501 vss 0.00786f
C3656 vdd.t275 vss 0.00385f
C3657 vdd.n63 vss 0.0167f
C3658 vdd.t417 vss 0.0098f
C3659 vdd.t378 vss 0.00522f
C3660 vdd.t439 vss 0.00522f
C3661 vdd.n64 vss 0.01114f
C3662 vdd.t376 vss 0.0198f
C3663 vdd.t274 vss 0.08979f
C3664 vdd.t500 vss 0.14646f
C3665 vdd.t416 vss 0.12034f
C3666 vdd.t499 vss 0.08209f
C3667 vdd.t415 vss 0.10355f
C3668 vdd.t438 vss 0.10355f
C3669 vdd.t377 vss 0.14739f
C3670 vdd.t375 vss 0.17025f
C3671 vdd.n65 vss 0.10679f
C3672 vdd.t394 vss 0.00786f
C3673 vdd.t522 vss 0.00385f
C3674 vdd.n66 vss 0.0167f
C3675 vdd.t398 vss 0.0098f
C3676 vdd.t136 vss 0.00522f
C3677 vdd.t129 vss 0.00522f
C3678 vdd.n67 vss 0.01114f
C3679 vdd.t138 vss 0.0198f
C3680 vdd.t431 vss 0.01707f
C3681 vdd.t511 vss 0.01684f
C3682 vdd.t503 vss 0.01948f
C3683 vdd.t521 vss 0.08979f
C3684 vdd.t393 vss 0.14646f
C3685 vdd.t397 vss 0.12034f
C3686 vdd.t392 vss 0.08209f
C3687 vdd.t57 vss 0.10355f
C3688 vdd.t128 vss 0.10355f
C3689 vdd.t135 vss 0.14739f
C3690 vdd.t137 vss 0.16115f
C3691 vdd.t430 vss 0.0723f
C3692 vdd.t510 vss 0.10588f
C3693 vdd.t502 vss 0.11495f
C3694 vdd.t408 vss 0.2944f
C3695 vdd.t327 vss 0.12528f
C3696 vdd.t298 vss 0.12528f
C3697 vdd.t344 vss 0.12528f
C3698 vdd.t296 vss 0.12528f
C3699 vdd.t329 vss 0.12528f
C3700 vdd.t346 vss 0.12528f
C3701 vdd.t343 vss 0.12528f
C3702 vdd.t326 vss 0.12528f
C3703 vdd.t297 vss 0.12528f
C3704 vdd.t211 vss 0.12528f
C3705 vdd.t325 vss 0.12528f
C3706 vdd.t210 vss 0.12528f
C3707 vdd.t345 vss 0.12528f
C3708 vdd.t324 vss 0.12528f
C3709 vdd.t498 vss 0.12528f
C3710 vdd.t295 vss 0.12528f
C3711 vdd.t328 vss 0.16571f
C3712 vdd.t25 vss 0.01948f
C3713 vdd.t24 vss 0.12758f
C3714 vdd.t350 vss 0.2944f
C3715 vdd.t420 vss 0.12528f
C3716 vdd.t422 vss 0.12528f
C3717 vdd.t351 vss 0.12528f
C3718 vdd.t529 vss 0.12528f
C3719 vdd.t358 vss 0.12528f
C3720 vdd.t479 vss 0.12528f
C3721 vdd.t433 vss 0.12528f
C3722 vdd.t310 vss 0.12528f
C3723 vdd.t421 vss 0.12528f
C3724 vdd.t342 vss 0.12528f
C3725 vdd.t311 vss 0.12528f
C3726 vdd.t530 vss 0.12528f
C3727 vdd.t359 vss 0.12528f
C3728 vdd.t480 vss 0.12528f
C3729 vdd.t291 vss 0.12528f
C3730 vdd.t118 vss 0.12528f
C3731 vdd.t432 vss 0.16571f
C3732 vdd.t400 vss 0.01948f
C3733 vdd.t399 vss 0.12758f
C3734 vdd.t466 vss 0.2944f
C3735 vdd.t464 vss 0.12528f
C3736 vdd.t477 vss 0.12528f
C3737 vdd.t43 vss 0.12528f
C3738 vdd.t465 vss 0.12528f
C3739 vdd.t478 vss 0.12528f
C3740 vdd.t531 vss 0.12528f
C3741 vdd.t486 vss 0.12528f
C3742 vdd.t20 vss 0.12528f
C3743 vdd.t467 vss 0.12528f
C3744 vdd.t19 vss 0.12528f
C3745 vdd.t463 vss 0.12528f
C3746 vdd.t468 vss 0.12528f
C3747 vdd.t484 vss 0.12528f
C3748 vdd.t532 vss 0.12528f
C3749 vdd.t17 vss 0.12528f
C3750 vdd.t18 vss 0.12528f
C3751 vdd.t485 vss 0.16571f
C3752 vdd.t241 vss 0.01948f
C3753 vdd.t240 vss 0.12758f
C3754 vdd.t84 vss 0.2944f
C3755 vdd.t77 vss 0.12528f
C3756 vdd.t73 vss 0.12528f
C3757 vdd.t81 vss 0.12528f
C3758 vdd.t74 vss 0.12528f
C3759 vdd.t71 vss 0.12528f
C3760 vdd.t80 vss 0.12528f
C3761 vdd.t79 vss 0.12528f
C3762 vdd.t70 vss 0.12528f
C3763 vdd.t68 vss 0.12528f
C3764 vdd.t83 vss 0.12528f
C3765 vdd.t76 vss 0.12528f
C3766 vdd.t72 vss 0.12528f
C3767 vdd.t82 vss 0.12528f
C3768 vdd.t75 vss 0.12528f
C3769 vdd.t78 vss 0.12528f
C3770 vdd.t69 vss 0.12528f
C3771 vdd.t85 vss 0.16571f
C3772 vdd.t46 vss 0.01948f
C3773 vdd.t45 vss 0.12758f
C3774 vdd.t259 vss 0.2944f
C3775 vdd.t218 vss 0.12528f
C3776 vdd.t215 vss 0.12528f
C3777 vdd.t260 vss 0.12528f
C3778 vdd.t237 vss 0.12528f
C3779 vdd.t221 vss 0.12528f
C3780 vdd.t252 vss 0.12528f
C3781 vdd.t258 vss 0.12528f
C3782 vdd.t222 vss 0.12528f
C3783 vdd.t253 vss 0.12528f
C3784 vdd.t217 vss 0.12528f
C3785 vdd.t208 vss 0.12528f
C3786 vdd.t219 vss 0.12528f
C3787 vdd.t207 vss 0.12528f
C3788 vdd.t388 vss 0.12528f
C3789 vdd.t220 vss 0.12528f
C3790 vdd.t251 vss 0.12528f
C3791 vdd.t216 vss 0.16571f
C3792 vdd.t64 vss 0.01948f
C3793 vdd.t63 vss 0.12758f
C3794 vdd.t276 vss 0.2944f
C3795 vdd.t225 vss 0.12528f
C3796 vdd.t61 vss 0.12528f
C3797 vdd.t277 vss 0.12528f
C3798 vdd.t332 vss 0.12528f
C3799 vdd.t236 vss 0.12528f
C3800 vdd.t10 vss 0.12528f
C3801 vdd.t539 vss 0.12528f
C3802 vdd.t227 vss 0.12528f
C3803 vdd.t60 vss 0.12528f
C3804 vdd.t62 vss 0.12528f
C3805 vdd.t228 vss 0.12528f
C3806 vdd.t235 vss 0.12528f
C3807 vdd.t8 vss 0.12528f
C3808 vdd.t537 vss 0.12528f
C3809 vdd.t226 vss 0.12528f
C3810 vdd.t9 vss 0.12528f
C3811 vdd.t538 vss 0.16571f
C3812 vdd.t22 vss 0.01948f
C3813 vdd.t21 vss 0.12758f
C3814 vdd.t206 vss 0.2944f
C3815 vdd.t213 vss 0.12528f
C3816 vdd.t248 vss 0.12528f
C3817 vdd.t361 vss 0.12528f
C3818 vdd.t205 vss 0.12528f
C3819 vdd.t249 vss 0.12528f
C3820 vdd.t362 vss 0.12528f
C3821 vdd.t202 vss 0.12528f
C3822 vdd.t154 vss 0.12528f
C3823 vdd.t214 vss 0.12528f
C3824 vdd.t360 vss 0.12528f
C3825 vdd.t212 vss 0.12528f
C3826 vdd.t247 vss 0.12528f
C3827 vdd.t198 vss 0.12528f
C3828 vdd.t200 vss 0.12528f
C3829 vdd.t250 vss 0.12528f
C3830 vdd.t199 vss 0.12528f
C3831 vdd.t201 vss 0.16571f
C3832 vdd.t497 vss 0.01948f
C3833 vdd.t496 vss 0.12758f
C3834 vdd.t352 vss 0.2944f
C3835 vdd.t302 vss 0.12528f
C3836 vdd.t209 vss 0.12528f
C3837 vdd.t491 vss 0.12528f
C3838 vdd.t333 vss 0.12528f
C3839 vdd.t507 vss 0.12528f
C3840 vdd.t187 vss 0.12528f
C3841 vdd.t334 vss 0.12528f
C3842 vdd.t292 vss 0.12528f
C3843 vdd.t238 vss 0.12528f
C3844 vdd.t162 vss 0.12528f
C3845 vdd.t163 vss 0.12528f
C3846 vdd.t239 vss 0.12528f
C3847 vdd.t278 vss 0.12528f
C3848 vdd.t403 vss 0.12528f
C3849 vdd.t353 vss 0.12528f
C3850 vdd.t303 vss 0.12528f
C3851 vdd.t188 vss 0.16571f
C3852 vdd.t108 vss 0.01948f
C3853 vdd.t107 vss 0.12758f
C3854 vdd.t349 vss 0.2944f
C3855 vdd.t308 vss 0.12528f
C3856 vdd.t341 vss 0.12528f
C3857 vdd.t300 vss 0.12528f
C3858 vdd.t337 vss 0.12528f
C3859 vdd.t355 vss 0.12528f
C3860 vdd.t357 vss 0.12528f
C3861 vdd.t348 vss 0.12528f
C3862 vdd.t299 vss 0.12528f
C3863 vdd.t261 vss 0.12528f
C3864 vdd.t488 vss 0.12528f
C3865 vdd.t301 vss 0.12528f
C3866 vdd.t338 vss 0.12528f
C3867 vdd.t356 vss 0.12528f
C3868 vdd.t347 vss 0.12528f
C3869 vdd.t354 vss 0.12528f
C3870 vdd.t309 vss 0.12528f
C3871 vdd.t487 vss 0.16571f
C3872 vdd.t396 vss 0.01948f
C3873 vdd.t395 vss 0.12758f
C3874 vdd.t505 vss 0.2944f
C3875 vdd.t204 vss 0.12528f
C3876 vdd.t314 vss 0.12528f
C3877 vdd.t506 vss 0.12528f
C3878 vdd.t401 vss 0.12528f
C3879 vdd.t330 vss 0.12528f
C3880 vdd.t312 vss 0.12528f
C3881 vdd.t391 vss 0.12528f
C3882 vdd.t245 vss 0.12528f
C3883 vdd.t313 vss 0.12528f
C3884 vdd.t504 vss 0.12528f
C3885 vdd.t203 vss 0.12528f
C3886 vdd.t402 vss 0.12528f
C3887 vdd.t331 vss 0.12528f
C3888 vdd.t389 vss 0.12528f
C3889 vdd.t244 vss 0.12528f
C3890 vdd.t246 vss 0.12528f
C3891 vdd.t390 vss 0.16571f
C3892 vdd.t230 vss 0.01948f
C3893 vdd.t229 vss 0.12758f
C3894 vdd.n68 vss 0.26018f
C3895 vdd.n69 vss 0.29969f
C3896 vdd.n70 vss 0.51554f
C3897 vdd.n71 vss 0.2591f
C3898 vdd.n72 vss 0.28357f
C3899 vdd.n73 vss 0.49515f
C3900 vdd.n74 vss 0.2591f
C3901 vdd.n75 vss 0.28357f
C3902 vdd.n76 vss 0.49515f
C3903 vdd.n77 vss 0.2591f
C3904 vdd.n78 vss 0.28357f
C3905 vdd.n79 vss 0.49515f
C3906 vdd.n80 vss 0.2591f
C3907 vdd.n81 vss 0.28357f
C3908 vdd.n82 vss 0.49515f
C3909 vdd.n83 vss 0.2591f
C3910 vdd.n84 vss 0.28357f
C3911 vdd.n85 vss 0.49515f
C3912 vdd.n86 vss 0.2591f
C3913 vdd.n87 vss 0.28357f
C3914 vdd.n88 vss 0.49515f
C3915 vdd.n89 vss 0.2591f
C3916 vdd.n90 vss 0.28357f
C3917 vdd.n91 vss 0.49515f
C3918 vdd.n92 vss 0.2591f
C3919 vdd.n93 vss 0.28357f
C3920 vdd.n94 vss 0.49515f
C3921 vdd.n95 vss 0.2591f
C3922 vdd.n96 vss 0.28357f
C3923 vdd.n97 vss 0.62307f
C3924 vdd.n98 vss 0.3655f
C3925 vdd.n99 vss 0.05225f
C3926 vdd.n100 vss 0.04503f
C3927 vdd.n101 vss 0.04754f
C3928 vdd.n102 vss 0.06466f
C3929 vdd.n103 vss 0.10166f
C3930 vdd.n104 vss 0.09174f
C3931 vdd.n105 vss 0.06315f
C3932 vdd.n106 vss 0.05676f
C3933 vdd.n107 vss 0.06669f
C3934 vdd.n108 vss 0.10166f
C3935 vdd.n109 vss 0.09174f
C3936 vdd.n110 vss 0.04468f
C3937 vdd.n111 vss 0.04524f
C3938 vdd.n112 vss 0.05663f
C3939 vdd.n113 vss 0.05225f
C3940 vdd.n114 vss 0.04503f
C3941 vdd.n115 vss 0.04754f
C3942 vdd.n116 vss 0.06466f
C3943 vdd.n117 vss 0.10166f
C3944 vdd.n118 vss 0.09174f
C3945 vdd.n119 vss 0.06315f
C3946 vdd.n120 vss 0.05676f
C3947 vdd.n121 vss 0.06669f
C3948 vdd.n122 vss 0.10166f
C3949 vdd.n123 vss 0.09174f
C3950 vdd.n124 vss 0.04468f
C3951 vdd.n125 vss 0.04524f
C3952 vdd.n126 vss 0.05663f
C3953 vdd.n127 vss 0.05225f
C3954 vdd.n128 vss 0.04503f
C3955 vdd.n129 vss 0.04754f
C3956 vdd.n130 vss 0.06466f
C3957 vdd.n131 vss 0.10166f
C3958 vdd.n132 vss 0.09174f
C3959 vdd.n133 vss 0.06315f
C3960 vdd.n134 vss 0.05676f
C3961 vdd.n135 vss 0.06669f
C3962 vdd.n136 vss 0.10166f
C3963 vdd.n137 vss 0.09174f
C3964 vdd.n138 vss 0.04468f
C3965 vdd.n139 vss 0.04524f
C3966 vdd.n140 vss 0.05663f
C3967 vdd.n141 vss 0.05225f
C3968 vdd.n142 vss 0.04503f
C3969 vdd.n143 vss 0.04754f
C3970 vdd.n144 vss 0.06466f
C3971 vdd.n145 vss 0.10166f
C3972 vdd.n146 vss 0.09174f
C3973 vdd.n147 vss 0.06315f
C3974 vdd.n148 vss 0.05676f
C3975 vdd.n149 vss 0.06669f
C3976 vdd.n150 vss 0.10166f
C3977 vdd.n151 vss 0.09174f
C3978 vdd.n152 vss 0.04468f
C3979 vdd.n153 vss 0.04524f
C3980 vdd.n154 vss 0.05663f
C3981 vdd.n155 vss 0.05225f
C3982 vdd.n156 vss 0.04503f
C3983 vdd.n157 vss 0.04754f
C3984 vdd.n158 vss 0.06466f
C3985 vdd.n159 vss 0.10166f
C3986 vdd.n160 vss 0.09174f
C3987 vdd.n161 vss 0.06315f
C3988 vdd.n162 vss 0.05676f
C3989 vdd.n163 vss 0.06669f
C3990 vdd.n164 vss 0.10166f
C3991 vdd.n165 vss 0.09174f
C3992 vdd.n166 vss 0.04468f
C3993 vdd.n167 vss 0.04524f
C3994 vdd.n168 vss 0.05663f
C3995 vdd.n169 vss 0.05225f
C3996 vdd.n170 vss 0.04503f
C3997 vdd.n171 vss 0.04754f
C3998 vdd.n172 vss 0.06466f
C3999 vdd.n173 vss 0.10166f
C4000 vdd.n174 vss 0.09174f
C4001 vdd.n175 vss 0.06315f
C4002 vdd.n176 vss 0.05676f
C4003 vdd.n177 vss 0.06669f
C4004 vdd.n178 vss 0.10166f
C4005 vdd.n179 vss 0.09174f
C4006 vdd.n180 vss 0.04468f
C4007 vdd.n181 vss 0.04524f
C4008 vdd.n182 vss 0.05663f
C4009 vdd.n183 vss 0.05225f
C4010 vdd.n184 vss 0.04503f
C4011 vdd.n185 vss 0.04754f
C4012 vdd.n186 vss 0.06466f
C4013 vdd.n187 vss 0.10166f
C4014 vdd.n188 vss 0.09174f
C4015 vdd.n189 vss 0.06315f
C4016 vdd.n190 vss 0.05676f
C4017 vdd.n191 vss 0.06669f
C4018 vdd.n192 vss 0.10166f
C4019 vdd.n193 vss 0.09174f
C4020 vdd.n194 vss 0.04468f
C4021 vdd.n195 vss 0.04524f
C4022 vdd.n196 vss 0.05663f
C4023 vdd.n197 vss 0.05225f
C4024 vdd.n198 vss 0.04503f
C4025 vdd.n199 vss 0.04754f
C4026 vdd.n200 vss 0.06466f
C4027 vdd.n201 vss 0.10166f
C4028 vdd.n202 vss 0.09174f
C4029 vdd.n203 vss 0.06315f
C4030 vdd.n204 vss 0.05676f
C4031 vdd.n205 vss 0.06669f
C4032 vdd.n206 vss 0.10166f
C4033 vdd.n207 vss 0.09174f
C4034 vdd.n208 vss 0.04468f
C4035 vdd.n209 vss 0.04524f
C4036 vdd.n210 vss 0.05663f
C4037 vdd.n211 vss 0.05225f
C4038 vdd.n212 vss 0.04503f
C4039 vdd.n213 vss 0.04754f
C4040 vdd.n214 vss 0.06466f
C4041 vdd.n215 vss 0.10166f
C4042 vdd.n216 vss 0.09174f
C4043 vdd.n217 vss 0.06315f
C4044 vdd.n218 vss 0.05676f
C4045 vdd.n219 vss 0.06669f
C4046 vdd.n220 vss 0.10166f
C4047 vdd.n221 vss 0.09174f
C4048 vdd.n222 vss 0.04468f
C4049 vdd.n223 vss 0.04524f
C4050 vdd.n224 vss 0.05663f
C4051 vdd.n225 vss 0.05225f
C4052 vdd.n226 vss 0.04503f
C4053 vdd.n227 vss 0.04754f
C4054 vdd.n228 vss 0.06466f
C4055 vdd.n229 vss 0.10166f
C4056 vdd.n230 vss 0.09174f
C4057 vdd.n231 vss 0.06315f
C4058 vdd.n232 vss 0.05676f
C4059 vdd.n233 vss 0.06669f
C4060 vdd.n234 vss 0.10166f
C4061 vdd.n235 vss 0.09174f
C4062 vdd.n236 vss 0.04468f
C4063 vdd.n237 vss 0.17012f
C4064 pin.t96 vss 0.52415f
C4065 pin.t99 vss 0.07403f
C4066 pin.t95 vss 0.07403f
C4067 pin.n0 vss 0.34895f
C4068 pin.t94 vss 0.07403f
C4069 pin.t97 vss 0.07403f
C4070 pin.n1 vss 0.34895f
C4071 pin.t98 vss 0.52415f
C4072 pin.t230 vss 0.54448f
C4073 pin.t145 vss 0.07403f
C4074 pin.t71 vss 0.07403f
C4075 pin.n2 vss 0.35196f
C4076 pin.t197 vss 0.07403f
C4077 pin.t231 vss 0.07403f
C4078 pin.n3 vss 0.35196f
C4079 pin.t143 vss 0.07403f
C4080 pin.t152 vss 0.07403f
C4081 pin.n4 vss 0.35196f
C4082 pin.t112 vss 0.07403f
C4083 pin.t184 vss 0.07403f
C4084 pin.n5 vss 0.35196f
C4085 pin.t229 vss 0.07403f
C4086 pin.t144 vss 0.07403f
C4087 pin.n6 vss 0.35196f
C4088 pin.t198 vss 0.07403f
C4089 pin.t70 vss 0.07403f
C4090 pin.n7 vss 0.35196f
C4091 pin.t182 vss 0.07403f
C4092 pin.t153 vss 0.07403f
C4093 pin.n8 vss 0.35196f
C4094 pin.t113 vss 0.07403f
C4095 pin.t111 vss 0.07403f
C4096 pin.n9 vss 0.35196f
C4097 pin.t183 vss 0.54448f
C4098 pin.t186 vss 0.52415f
C4099 pin.t189 vss 0.07403f
C4100 pin.t190 vss 0.07403f
C4101 pin.n10 vss 0.34895f
C4102 pin.t188 vss 0.07403f
C4103 pin.t185 vss 0.07403f
C4104 pin.n11 vss 0.34895f
C4105 pin.t187 vss 0.52415f
C4106 pin.t167 vss 0.54448f
C4107 pin.t159 vss 0.07403f
C4108 pin.t139 vss 0.07403f
C4109 pin.n12 vss 0.35196f
C4110 pin.t157 vss 0.07403f
C4111 pin.t135 vss 0.07403f
C4112 pin.n13 vss 0.35196f
C4113 pin.t175 vss 0.07403f
C4114 pin.t173 vss 0.07403f
C4115 pin.n14 vss 0.35196f
C4116 pin.t134 vss 0.07403f
C4117 pin.t166 vss 0.07403f
C4118 pin.n15 vss 0.35196f
C4119 pin.t220 vss 0.07403f
C4120 pin.t124 vss 0.07403f
C4121 pin.n16 vss 0.35196f
C4122 pin.t158 vss 0.07403f
C4123 pin.t136 vss 0.07403f
C4124 pin.n17 vss 0.35196f
C4125 pin.t165 vss 0.07403f
C4126 pin.t174 vss 0.07403f
C4127 pin.n18 vss 0.35196f
C4128 pin.t140 vss 0.07403f
C4129 pin.t172 vss 0.07403f
C4130 pin.n19 vss 0.35196f
C4131 pin.t219 vss 0.54448f
C4132 pin.t57 vss 0.52415f
C4133 pin.t53 vss 0.07403f
C4134 pin.t54 vss 0.07403f
C4135 pin.n20 vss 0.34895f
C4136 pin.t58 vss 0.07403f
C4137 pin.t56 vss 0.07403f
C4138 pin.n21 vss 0.34895f
C4139 pin.t55 vss 0.52415f
C4140 pin.t170 vss 0.54448f
C4141 pin.t76 vss 0.07403f
C4142 pin.t137 vss 0.07403f
C4143 pin.n22 vss 0.35196f
C4144 pin.t155 vss 0.07403f
C4145 pin.t221 vss 0.07403f
C4146 pin.n23 vss 0.35196f
C4147 pin.t63 vss 0.07403f
C4148 pin.t232 vss 0.07403f
C4149 pin.n24 vss 0.35196f
C4150 pin.t129 vss 0.07403f
C4151 pin.t156 vss 0.07403f
C4152 pin.n25 vss 0.35196f
C4153 pin.t61 vss 0.07403f
C4154 pin.t103 vss 0.07403f
C4155 pin.n26 vss 0.35196f
C4156 pin.t104 vss 0.07403f
C4157 pin.t62 vss 0.07403f
C4158 pin.n27 vss 0.35196f
C4159 pin.t199 vss 0.07403f
C4160 pin.t127 vss 0.07403f
C4161 pin.n28 vss 0.35196f
C4162 pin.t138 vss 0.07403f
C4163 pin.t171 vss 0.07403f
C4164 pin.n29 vss 0.35196f
C4165 pin.t64 vss 0.54448f
C4166 pin.t226 vss 0.52415f
C4167 pin.t224 vss 0.07403f
C4168 pin.t223 vss 0.07403f
C4169 pin.n30 vss 0.34895f
C4170 pin.t222 vss 0.07403f
C4171 pin.t225 vss 0.07403f
C4172 pin.n31 vss 0.34895f
C4173 pin.t227 vss 0.52415f
C4174 pin.t73 vss 0.54448f
C4175 pin.t115 vss 0.07403f
C4176 pin.t80 vss 0.07403f
C4177 pin.n32 vss 0.35196f
C4178 pin.t72 vss 0.07403f
C4179 pin.t179 vss 0.07403f
C4180 pin.n33 vss 0.35196f
C4181 pin.t180 vss 0.07403f
C4182 pin.t116 vss 0.07403f
C4183 pin.n34 vss 0.35196f
C4184 pin.t60 vss 0.07403f
C4185 pin.t69 vss 0.07403f
C4186 pin.n35 vss 0.35196f
C4187 pin.t178 vss 0.07403f
C4188 pin.t81 vss 0.07403f
C4189 pin.n36 vss 0.35196f
C4190 pin.t114 vss 0.07403f
C4191 pin.t79 vss 0.07403f
C4192 pin.n37 vss 0.35196f
C4193 pin.t67 vss 0.07403f
C4194 pin.t65 vss 0.07403f
C4195 pin.n38 vss 0.35196f
C4196 pin.t66 vss 0.07403f
C4197 pin.t117 vss 0.07403f
C4198 pin.n39 vss 0.35196f
C4199 pin.t68 vss 0.54448f
C4200 pin.t10 vss 0.52415f
C4201 pin.t8 vss 0.07403f
C4202 pin.t12 vss 0.07403f
C4203 pin.n40 vss 0.34895f
C4204 pin.t9 vss 0.07403f
C4205 pin.t11 vss 0.07403f
C4206 pin.n41 vss 0.34895f
C4207 pin.t7 vss 0.52415f
C4208 pin.t125 vss 0.54448f
C4209 pin.t27 vss 0.07403f
C4210 pin.t90 vss 0.07403f
C4211 pin.n42 vss 0.35196f
C4212 pin.t154 vss 0.07403f
C4213 pin.t126 vss 0.07403f
C4214 pin.n43 vss 0.35196f
C4215 pin.t2 vss 0.07403f
C4216 pin.t101 vss 0.07403f
C4217 pin.n44 vss 0.35196f
C4218 pin.t92 vss 0.07403f
C4219 pin.t239 vss 0.07403f
C4220 pin.n45 vss 0.35196f
C4221 pin.t28 vss 0.07403f
C4222 pin.t26 vss 0.07403f
C4223 pin.n46 vss 0.35196f
C4224 pin.t100 vss 0.07403f
C4225 pin.t93 vss 0.07403f
C4226 pin.n47 vss 0.35196f
C4227 pin.t237 vss 0.07403f
C4228 pin.t0 vss 0.07403f
C4229 pin.n48 vss 0.35196f
C4230 pin.t1 vss 0.07403f
C4231 pin.t91 vss 0.07403f
C4232 pin.n49 vss 0.35196f
C4233 pin.t238 vss 0.54448f
C4234 pin.t31 vss 0.52415f
C4235 pin.t34 vss 0.07403f
C4236 pin.t30 vss 0.07403f
C4237 pin.n50 vss 0.34895f
C4238 pin.t29 vss 0.07403f
C4239 pin.t32 vss 0.07403f
C4240 pin.n51 vss 0.34895f
C4241 pin.t33 vss 0.52415f
C4242 pin.t122 vss 0.54448f
C4243 pin.t82 vss 0.07403f
C4244 pin.t85 vss 0.07403f
C4245 pin.n52 vss 0.35196f
C4246 pin.t102 vss 0.07403f
C4247 pin.t123 vss 0.07403f
C4248 pin.n53 vss 0.35196f
C4249 pin.t119 vss 0.07403f
C4250 pin.t88 vss 0.07403f
C4251 pin.n54 vss 0.35196f
C4252 pin.t89 vss 0.07403f
C4253 pin.t121 vss 0.07403f
C4254 pin.n55 vss 0.35196f
C4255 pin.t84 vss 0.07403f
C4256 pin.t120 vss 0.07403f
C4257 pin.n56 vss 0.35196f
C4258 pin.t86 vss 0.07403f
C4259 pin.t75 vss 0.07403f
C4260 pin.n57 vss 0.35196f
C4261 pin.t181 vss 0.07403f
C4262 pin.t74 vss 0.07403f
C4263 pin.n58 vss 0.35196f
C4264 pin.t118 vss 0.07403f
C4265 pin.t87 vss 0.07403f
C4266 pin.n59 vss 0.35196f
C4267 pin.t83 vss 0.54448f
C4268 pin.t21 vss 0.52415f
C4269 pin.t22 vss 0.07403f
C4270 pin.t23 vss 0.07403f
C4271 pin.n60 vss 0.34895f
C4272 pin.t25 vss 0.07403f
C4273 pin.t20 vss 0.07403f
C4274 pin.n61 vss 0.34895f
C4275 pin.t24 vss 0.52415f
C4276 pin.t51 vss 0.54448f
C4277 pin.t40 vss 0.07403f
C4278 pin.t44 vss 0.07403f
C4279 pin.n62 vss 0.35196f
C4280 pin.t41 vss 0.07403f
C4281 pin.t48 vss 0.07403f
C4282 pin.n63 vss 0.35196f
C4283 pin.t47 vss 0.07403f
C4284 pin.t38 vss 0.07403f
C4285 pin.n64 vss 0.35196f
C4286 pin.t37 vss 0.07403f
C4287 pin.t46 vss 0.07403f
C4288 pin.n65 vss 0.35196f
C4289 pin.t50 vss 0.07403f
C4290 pin.t35 vss 0.07403f
C4291 pin.n66 vss 0.35196f
C4292 pin.t39 vss 0.07403f
C4293 pin.t43 vss 0.07403f
C4294 pin.n67 vss 0.35196f
C4295 pin.t42 vss 0.07403f
C4296 pin.t49 vss 0.07403f
C4297 pin.n68 vss 0.35196f
C4298 pin.t36 vss 0.07403f
C4299 pin.t45 vss 0.07403f
C4300 pin.n69 vss 0.35196f
C4301 pin.t52 vss 0.54448f
C4302 pin.t106 vss 0.52415f
C4303 pin.t107 vss 0.07403f
C4304 pin.t108 vss 0.07403f
C4305 pin.n70 vss 0.34895f
C4306 pin.t110 vss 0.07403f
C4307 pin.t105 vss 0.07403f
C4308 pin.n71 vss 0.34895f
C4309 pin.t109 vss 0.52415f
C4310 pin.t209 vss 0.54448f
C4311 pin.t212 vss 0.07403f
C4312 pin.t207 vss 0.07403f
C4313 pin.n72 vss 0.35196f
C4314 pin.t208 vss 0.07403f
C4315 pin.t19 vss 0.07403f
C4316 pin.n73 vss 0.35196f
C4317 pin.t235 vss 0.07403f
C4318 pin.t213 vss 0.07403f
C4319 pin.n74 vss 0.35196f
C4320 pin.t6 vss 0.07403f
C4321 pin.t218 vss 0.07403f
C4322 pin.n75 vss 0.35196f
C4323 pin.t5 vss 0.07403f
C4324 pin.t210 vss 0.07403f
C4325 pin.n76 vss 0.35196f
C4326 pin.t211 vss 0.07403f
C4327 pin.t206 vss 0.07403f
C4328 pin.n77 vss 0.35196f
C4329 pin.t236 vss 0.07403f
C4330 pin.t216 vss 0.07403f
C4331 pin.n78 vss 0.35196f
C4332 pin.t4 vss 0.07403f
C4333 pin.t3 vss 0.07403f
C4334 pin.n79 vss 0.35196f
C4335 pin.t217 vss 0.54448f
C4336 pin.t192 vss 0.52415f
C4337 pin.t196 vss 0.07403f
C4338 pin.t191 vss 0.07403f
C4339 pin.n80 vss 0.34895f
C4340 pin.t193 vss 0.07403f
C4341 pin.t194 vss 0.07403f
C4342 pin.n81 vss 0.34895f
C4343 pin.t195 vss 0.52415f
C4344 pin.t168 vss 0.54448f
C4345 pin.t203 vss 0.07403f
C4346 pin.t201 vss 0.07403f
C4347 pin.n82 vss 0.35196f
C4348 pin.t233 vss 0.07403f
C4349 pin.t169 vss 0.07403f
C4350 pin.n83 vss 0.35196f
C4351 pin.t214 vss 0.07403f
C4352 pin.t176 vss 0.07403f
C4353 pin.n84 vss 0.35196f
C4354 pin.t141 vss 0.07403f
C4355 pin.t205 vss 0.07403f
C4356 pin.n85 vss 0.35196f
C4357 pin.t160 vss 0.07403f
C4358 pin.t202 vss 0.07403f
C4359 pin.n86 vss 0.35196f
C4360 pin.t234 vss 0.07403f
C4361 pin.t142 vss 0.07403f
C4362 pin.n87 vss 0.35196f
C4363 pin.t215 vss 0.07403f
C4364 pin.t177 vss 0.07403f
C4365 pin.n88 vss 0.35196f
C4366 pin.t59 vss 0.07403f
C4367 pin.t128 vss 0.07403f
C4368 pin.n89 vss 0.35196f
C4369 pin.t204 vss 0.54448f
C4370 pin.t15 vss 0.52415f
C4371 pin.t14 vss 0.07403f
C4372 pin.t18 vss 0.07403f
C4373 pin.n90 vss 0.34895f
C4374 pin.t17 vss 0.07403f
C4375 pin.t16 vss 0.07403f
C4376 pin.n91 vss 0.34895f
C4377 pin.t13 vss 0.52415f
C4378 pin.t200 vss 0.54448f
C4379 pin.t133 vss 0.07403f
C4380 pin.t149 vss 0.07403f
C4381 pin.n92 vss 0.35196f
C4382 pin.t131 vss 0.07403f
C4383 pin.t162 vss 0.07403f
C4384 pin.n93 vss 0.35196f
C4385 pin.t164 vss 0.07403f
C4386 pin.t151 vss 0.07403f
C4387 pin.n94 vss 0.35196f
C4388 pin.t148 vss 0.07403f
C4389 pin.t161 vss 0.07403f
C4390 pin.n95 vss 0.35196f
C4391 pin.t78 vss 0.07403f
C4392 pin.t132 vss 0.07403f
C4393 pin.n96 vss 0.35196f
C4394 pin.t77 vss 0.07403f
C4395 pin.t147 vss 0.07403f
C4396 pin.n97 vss 0.35196f
C4397 pin.t146 vss 0.07403f
C4398 pin.t163 vss 0.07403f
C4399 pin.n98 vss 0.35196f
C4400 pin.t130 vss 0.07403f
C4401 pin.t228 vss 0.07403f
C4402 pin.n99 vss 0.35196f
C4403 pin.t150 vss 0.55911f
C4404 pin.n100 vss 1.01244f
C4405 pin.n101 vss 0.28662f
C4406 pin.n102 vss 0.28662f
C4407 pin.n103 vss 0.28662f
C4408 pin.n104 vss 0.28662f
C4409 pin.n105 vss 0.28662f
C4410 pin.n106 vss 0.28662f
C4411 pin.n107 vss 0.29394f
C4412 pin.n108 vss 0.34424f
C4413 pin.n109 vss 0.34126f
C4414 pin.n110 vss 0.29641f
C4415 pin.n111 vss 0.29568f
C4416 pin.n112 vss 0.45122f
C4417 pin.n113 vss 0.49443f
C4418 pin.n114 vss 0.29394f
C4419 pin.n115 vss 0.28662f
C4420 pin.n116 vss 0.28662f
C4421 pin.n117 vss 0.28662f
C4422 pin.n118 vss 0.28662f
C4423 pin.n119 vss 0.28662f
C4424 pin.n120 vss 0.28662f
C4425 pin.n121 vss 0.29394f
C4426 pin.n122 vss 0.34424f
C4427 pin.n123 vss 0.34126f
C4428 pin.n124 vss 0.29641f
C4429 pin.n125 vss 0.29568f
C4430 pin.n126 vss 0.45122f
C4431 pin.n127 vss 0.49443f
C4432 pin.n128 vss 0.29394f
C4433 pin.n129 vss 0.28662f
C4434 pin.n130 vss 0.28662f
C4435 pin.n131 vss 0.28662f
C4436 pin.n132 vss 0.28662f
C4437 pin.n133 vss 0.28662f
C4438 pin.n134 vss 0.28662f
C4439 pin.n135 vss 0.29394f
C4440 pin.n136 vss 0.34424f
C4441 pin.n137 vss 0.34126f
C4442 pin.n138 vss 0.29641f
C4443 pin.n139 vss 0.29568f
C4444 pin.n140 vss 0.45122f
C4445 pin.n141 vss 0.49443f
C4446 pin.n142 vss 0.29394f
C4447 pin.n143 vss 0.28662f
C4448 pin.n144 vss 0.28662f
C4449 pin.n145 vss 0.28662f
C4450 pin.n146 vss 0.28662f
C4451 pin.n147 vss 0.28662f
C4452 pin.n148 vss 0.28662f
C4453 pin.n149 vss 0.29394f
C4454 pin.n150 vss 0.34424f
C4455 pin.n151 vss 0.34126f
C4456 pin.n152 vss 0.29641f
C4457 pin.n153 vss 0.29568f
C4458 pin.n154 vss 0.45122f
C4459 pin.n155 vss 0.49443f
C4460 pin.n156 vss 0.29394f
C4461 pin.n157 vss 0.28662f
C4462 pin.n158 vss 0.28662f
C4463 pin.n159 vss 0.28662f
C4464 pin.n160 vss 0.28662f
C4465 pin.n161 vss 0.28662f
C4466 pin.n162 vss 0.28662f
C4467 pin.n163 vss 0.29394f
C4468 pin.n164 vss 0.34424f
C4469 pin.n165 vss 0.34126f
C4470 pin.n166 vss 0.29641f
C4471 pin.n167 vss 0.29568f
C4472 pin.n168 vss 0.45122f
C4473 pin.n169 vss 0.49443f
C4474 pin.n170 vss 0.29394f
C4475 pin.n171 vss 0.28662f
C4476 pin.n172 vss 0.28662f
C4477 pin.n173 vss 0.28662f
C4478 pin.n174 vss 0.28662f
C4479 pin.n175 vss 0.28662f
C4480 pin.n176 vss 0.28662f
C4481 pin.n177 vss 0.29394f
C4482 pin.n178 vss 0.34424f
C4483 pin.n179 vss 0.34126f
C4484 pin.n180 vss 0.29641f
C4485 pin.n181 vss 0.29568f
C4486 pin.n182 vss 0.45122f
C4487 pin.n183 vss 0.49443f
C4488 pin.n184 vss 0.29394f
C4489 pin.n185 vss 0.28662f
C4490 pin.n186 vss 0.28662f
C4491 pin.n187 vss 0.28662f
C4492 pin.n188 vss 0.28662f
C4493 pin.n189 vss 0.28662f
C4494 pin.n190 vss 0.28662f
C4495 pin.n191 vss 0.29394f
C4496 pin.n192 vss 0.34424f
C4497 pin.n193 vss 0.34126f
C4498 pin.n194 vss 0.29641f
C4499 pin.n195 vss 0.29568f
C4500 pin.n196 vss 0.45122f
C4501 pin.n197 vss 0.49443f
C4502 pin.n198 vss 0.29394f
C4503 pin.n199 vss 0.28662f
C4504 pin.n200 vss 0.28662f
C4505 pin.n201 vss 0.28662f
C4506 pin.n202 vss 0.28662f
C4507 pin.n203 vss 0.28662f
C4508 pin.n204 vss 0.28662f
C4509 pin.n205 vss 0.29394f
C4510 pin.n206 vss 0.34424f
C4511 pin.n207 vss 0.34126f
C4512 pin.n208 vss 0.29641f
C4513 pin.n209 vss 0.29568f
C4514 pin.n210 vss 0.45122f
C4515 pin.n211 vss 0.49443f
C4516 pin.n212 vss 0.29394f
C4517 pin.n213 vss 0.28662f
C4518 pin.n214 vss 0.28662f
C4519 pin.n215 vss 0.28662f
C4520 pin.n216 vss 0.28662f
C4521 pin.n217 vss 0.28662f
C4522 pin.n218 vss 0.28662f
C4523 pin.n219 vss 0.29394f
C4524 pin.n220 vss 0.34424f
C4525 pin.n221 vss 0.34126f
C4526 pin.n222 vss 0.29641f
C4527 pin.n223 vss 0.29568f
C4528 pin.n224 vss 0.45122f
C4529 pin.n225 vss 0.57456f
C4530 pin.n226 vss 0.29394f
C4531 pin.n227 vss 0.28662f
C4532 pin.n228 vss 0.28662f
C4533 pin.n229 vss 0.28662f
C4534 pin.n230 vss 0.28662f
C4535 pin.n231 vss 0.28662f
C4536 pin.n232 vss 0.28662f
C4537 pin.n233 vss 0.29394f
C4538 pin.n234 vss 0.34424f
C4539 pin.n235 vss 0.34126f
C4540 pin.n236 vss 0.29641f
C4541 pin.n237 vss 0.29568f
C4542 pin.n238 vss 0.45122f
C4543 BUS[7].t3 vss 0.08734f
C4544 BUS[7].t1 vss 0.08734f
C4545 BUS[7].n0 vss 0.4704f
C4546 BUS[7].t0 vss 0.08734f
C4547 BUS[7].t2 vss 0.08734f
C4548 BUS[7].n1 vss 0.46764f
C4549 BUS[7].n2 vss 0.27386f
C4550 BUS[7].t4 vss 0.08734f
C4551 BUS[7].t5 vss 0.08734f
C4552 BUS[7].n3 vss 0.46764f
C4553 BUS[7].n4 vss 0.23641f
C4554 BUS[7].t18 vss 0.08734f
C4555 BUS[7].t15 vss 0.08734f
C4556 BUS[7].n5 vss 0.47045f
C4557 BUS[7].n6 vss 0.20977f
C4558 BUS[7].t16 vss 0.08734f
C4559 BUS[7].t6 vss 0.08734f
C4560 BUS[7].n7 vss 0.47317f
C4561 BUS[7].t19 vss 0.08734f
C4562 BUS[7].t12 vss 0.08734f
C4563 BUS[7].n8 vss 0.47045f
C4564 BUS[7].n9 vss 0.26765f
C4565 BUS[7].t23 vss 0.08734f
C4566 BUS[7].t9 vss 0.08734f
C4567 BUS[7].n10 vss 0.47045f
C4568 BUS[7].n11 vss 0.15534f
C4569 BUS[7].t17 vss 0.08734f
C4570 BUS[7].t14 vss 0.08734f
C4571 BUS[7].n12 vss 0.47045f
C4572 BUS[7].n13 vss 0.15534f
C4573 BUS[7].t13 vss 0.08734f
C4574 BUS[7].t7 vss 0.08734f
C4575 BUS[7].n14 vss 0.47045f
C4576 BUS[7].n15 vss 0.15534f
C4577 BUS[7].t20 vss 0.08734f
C4578 BUS[7].t21 vss 0.08734f
C4579 BUS[7].n16 vss 0.47045f
C4580 BUS[7].n17 vss 0.15534f
C4581 BUS[7].t8 vss 0.08734f
C4582 BUS[7].t11 vss 0.08734f
C4583 BUS[7].n18 vss 0.47045f
C4584 BUS[7].n19 vss 0.15534f
C4585 BUS[7].t22 vss 0.08734f
C4586 BUS[7].t10 vss 0.08734f
C4587 BUS[7].n20 vss 0.47045f
C4588 BUS[7].n21 vss 0.10378f
C4589 BUS[7].n22 vss 0.3948f
C4590 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t1 vss 0.06869f
C4591 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t0 vss 0.09485f
C4592 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t2 vss 0.12308f
C4593 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t18 vss 0.12285f
C4594 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n0 vss 0.18852f
C4595 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t9 vss 0.12285f
C4596 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n1 vss 0.10017f
C4597 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t12 vss 0.12285f
C4598 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n2 vss 0.10017f
C4599 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t5 vss 0.12285f
C4600 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n3 vss 0.10017f
C4601 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t15 vss 0.12285f
C4602 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n4 vss 0.10017f
C4603 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t11 vss 0.12285f
C4604 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n5 vss 0.10017f
C4605 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t4 vss 0.12285f
C4606 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n6 vss 0.10017f
C4607 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t19 vss 0.12285f
C4608 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n7 vss 0.10017f
C4609 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t17 vss 0.12285f
C4610 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n8 vss 0.10017f
C4611 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t8 vss 0.12285f
C4612 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n9 vss 0.10017f
C4613 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t7 vss 0.12285f
C4614 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n10 vss 0.10017f
C4615 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t16 vss 0.12285f
C4616 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n11 vss 0.10017f
C4617 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t13 vss 0.12285f
C4618 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n12 vss 0.10017f
C4619 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t6 vss 0.12285f
C4620 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n13 vss 0.10017f
C4621 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t14 vss 0.12285f
C4622 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n14 vss 0.10017f
C4623 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t10 vss 0.12285f
C4624 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n15 vss 0.10017f
C4625 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.t3 vss 0.12285f
C4626 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n16 vss 0.47233f
C4627 swmatrix_Tgate_0.gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0.ZN.n17 vss 0.46794f
.ends

