** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_row_10/swmatrix_row_10.sch
.subckt swmatrix_row_10 D_out D_in PHI_1 PHI_2 enable BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] VDD
+ pin VSS
*.PININFO pin:B PHI_2:I PHI_1:I BUS[1:10]:B D_in:I D_out:O VDD:B VSS:B enable:I
xSR D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] D_out gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8] gc[9] gc[10] PHI_1
+ PHI_2 enable VDD VSS ShiftReg_row_10_2
xTgates[1] gc[1] BUS[1] pin VSS VDD swmatrix_Tgate
xTgates[2] gc[2] BUS[2] pin VSS VDD swmatrix_Tgate
xTgates[3] gc[3] BUS[3] pin VSS VDD swmatrix_Tgate
xTgates[4] gc[4] BUS[4] pin VSS VDD swmatrix_Tgate
xTgates[5] gc[5] BUS[5] pin VSS VDD swmatrix_Tgate
xTgates[6] gc[6] BUS[6] pin VSS VDD swmatrix_Tgate
xTgates[7] gc[7] BUS[7] pin VSS VDD swmatrix_Tgate
xTgates[8] gc[8] BUS[8] pin VSS VDD swmatrix_Tgate
xTgates[9] gc[9] BUS[9] pin VSS VDD swmatrix_Tgate
xTgates[10] gc[10] BUS[10] pin VSS VDD swmatrix_Tgate
.ends

* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sch
.subckt ShiftReg_row_10_2 D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8]
+ gc[9] gc[10] PHI_1 PHI_2 EN VDD VSS
*.PININFO PHI_1:I PHI_2:I D_in:I Q[1:10]:O VDD:B VSS:B EN:B gc[1:10]:B
xFF[1] Q[1] D_in PHI_1 gc[1] PHI_2 EN VDD VSS DFF_2phase_1
xFF[2] Q[2] Q[1] PHI_1 gc[2] PHI_2 EN VDD VSS DFF_2phase_1
xFF[3] Q[3] Q[2] PHI_1 gc[3] PHI_2 EN VDD VSS DFF_2phase_1
xFF[4] Q[4] Q[3] PHI_1 gc[4] PHI_2 EN VDD VSS DFF_2phase_1
xFF[5] Q[5] Q[4] PHI_1 gc[5] PHI_2 EN VDD VSS DFF_2phase_1
xFF[6] Q[6] Q[5] PHI_1 gc[6] PHI_2 EN VDD VSS DFF_2phase_1
xFF[7] Q[7] Q[6] PHI_1 gc[7] PHI_2 EN VDD VSS DFF_2phase_1
xFF[8] Q[8] Q[7] PHI_1 gc[8] PHI_2 EN VDD VSS DFF_2phase_1
xFF[9] Q[9] Q[8] PHI_1 gc[9] PHI_2 EN VDD VSS DFF_2phase_1
xFF[10] Q[10] Q[9] PHI_1 gc[10] PHI_2 EN VDD VSS DFF_2phase_1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sym # of pins=5
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/swmatrix_Tgate/swmatrix_Tgate.sch
.subckt swmatrix_Tgate gated_control T2 T1 VSS VDD
*.PININFO T1:B T2:B VDD:B VSS:B gated_control:I
XM1 T1 gated_control T2 VSS nfet_03v3 L=0.28u W=24u nf=6 m=1
XM2 T1 gated_controlb T2 VDD pfet_03v3 L=0.28u W=68u nf=6 m=1
x1 gated_control gated_controlb VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends


* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 Q D PHI_1 gated_control PHI_2 EN VDD VSS
*.PININFO D:I PHI_1:I PHI_2:I Q:O VDD:B VSS:B gated_control:O EN:I
xmain D PHI_1 out_m VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
* noconn VSS
* noconn VDD
x1 net1 gated_control VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
x2 EN Q net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
.ends

