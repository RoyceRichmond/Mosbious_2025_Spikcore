** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/ShiftReg_row_10_2/ShiftReg_row_10_2.sch
.subckt DFF_10_row D_in Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8]
+ gc[9] gc[10] PHI_1 PHI_2 EN VDDd VSSd
*.PININFO PHI_1:I PHI_2:I D_in:I Q[1:10]:O VDDd:B VSSd:B EN:B gc[1:10]:B
xFF[1] Q[1] D_in PHI_1 gc[1] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[2] Q[2] Q[1] PHI_1 gc[2] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[3] Q[3] Q[2] PHI_1 gc[3] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[4] Q[4] Q[3] PHI_1 gc[4] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[5] Q[5] Q[4] PHI_1 gc[5] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[6] Q[6] Q[5] PHI_1 gc[6] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[7] Q[7] Q[6] PHI_1 gc[7] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[8] Q[8] Q[7] PHI_1 gc[8] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[9] Q[9] Q[8] PHI_1 gc[9] PHI_2 EN VDDd VSSd DFF_2phase_1
xFF[10] Q[10] Q[9] PHI_1 gc[10] PHI_2 EN VDDd VSSd DFF_2phase_1
.ends

* expanding   symbol:  designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym # of pins=8
** sym_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/Mosbious_2025_Spikcore/designs/libs/switch_matrix_gf180mcu_9t5v0/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 Q D PHI_1 gated_control PHI_2 EN VDDd VSSd
*.PININFO D:I PHI_1:I PHI_2:I Q:O VDDd:B VSSd:B gated_control:O EN:I
xmain D PHI_1 out_m VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
* noconn VSSd
* noconn VDDd
x1 net1 gated_control VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x2 EN Q net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
.ends

