* NGSPICE file created from swmatrix_row_10.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt DFF_2phase_1 gated_control PHI_1 D EN VDD Q PHI_2 VSS
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1_0 EN Q VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1_0/I
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q PHI_2 Q
+ VDD VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1$1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q
+ VDD VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1$1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0/I VDD VSS gated_control
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends

.subckt ShiftReg_row_10_2$1 VDD gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8] gc[9]
+ gc[10] Q[10] PHI_1 PHI_2 D_in Q[4] Q[9] Q[3] Q[8] Q[5] Q[7] Q[6] Q[1] Q[2] EN VSS
XDFF_2phase_1_0 gc[10] PHI_1 Q[9] EN VDD Q[10] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_1 gc[9] PHI_1 Q[8] EN VDD Q[9] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_2 gc[8] PHI_1 Q[7] EN VDD Q[8] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_3 gc[7] PHI_1 Q[6] EN VDD Q[7] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_4 gc[6] PHI_1 Q[5] EN VDD Q[6] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_5 gc[5] PHI_1 Q[4] EN VDD Q[5] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_6 gc[4] PHI_1 Q[3] EN VDD Q[4] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_7 gc[3] PHI_1 Q[2] EN VDD Q[3] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_8 gc[1] PHI_1 D_in EN VDD Q[1] PHI_2 VSS DFF_2phase_1
XDFF_2phase_1_9 gc[2] PHI_1 Q[1] EN VDD Q[2] PHI_2 VSS DFF_2phase_1
.ends

.subckt pfet a_1534_0# a_2174_0# a_1054_0# a_734_0# a_828_n136# a_28_n136# a_2588_n136#
+ a_1694_0# a_254_0# a_1628_n136# a_894_0# a_188_n136# a_988_n136# a_2814_0# a_2748_n136#
+ a_1788_n136# a_2334_0# a_348_n136# a_1214_0# a_1148_n136# a_1854_0# a_414_0# a_2108_n136#
+ a_2494_0# a_n92_0# a_1948_n136# a_1374_0# a_94_0# a_574_0# a_508_n136# a_2268_n136#
+ a_1308_n136# a_2014_0# a_668_n136# a_2428_n136# a_1468_n136# a_2654_0# w_n230_n138#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1 a_2654_0# a_2588_n136# a_2494_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X2 a_734_0# a_668_n136# a_574_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X3 a_2494_0# a_2428_n136# a_2334_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X4 a_254_0# a_188_n136# a_94_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X5 a_574_0# a_508_n136# a_414_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X6 a_2014_0# a_1948_n136# a_1854_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X7 a_1534_0# a_1468_n136# a_1374_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X8 a_1374_0# a_1308_n136# a_1214_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X9 a_1054_0# a_988_n136# a_894_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X10 a_2814_0# a_2748_n136# a_2654_0# w_n230_n138# pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X11 a_894_0# a_828_n136# a_734_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X12 a_2334_0# a_2268_n136# a_2174_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X13 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X14 a_2174_0# a_2108_n136# a_2014_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X15 a_414_0# a_348_n136# a_254_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X16 a_1854_0# a_1788_n136# a_1694_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X17 a_1694_0# a_1628_n136# a_1534_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt nfet vss a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_830_n132# a_414_0#
+ a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_350_n132#
X0 a_734_0# a_670_n132# a_574_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X3 a_894_0# a_830_n132# a_734_0# vss nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X4 a_94_0# a_30_n132# a_n84_0# vss nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X5 a_414_0# a_350_n132# a_254_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
.ends

.subckt swmatrix_Tgate VSS VDD T1 gated_control T2
Xpfet_0 T1 T1 T2 T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T2 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T1
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T1 T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ T1 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T2 T2 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN T2 VDD
+ pfet
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$1_0 gated_control VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$1
Xnfet_0 VSS T2 gated_control T1 T1 gated_control gated_control T2 gated_control T1
+ T2 gated_control T1 gated_control nfet
.ends

.subckt swmatrix_row_10 pin BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] d_out
XShiftReg_row_10_2$1_0 swmatrix_Tgate_9/VDD ShiftReg_row_10_2$1_0/gc[1] ShiftReg_row_10_2$1_0/gc[2]
+ ShiftReg_row_10_2$1_0/gc[3] ShiftReg_row_10_2$1_0/gc[4] ShiftReg_row_10_2$1_0/gc[5]
+ ShiftReg_row_10_2$1_0/gc[6] ShiftReg_row_10_2$1_0/gc[7] ShiftReg_row_10_2$1_0/gc[8]
+ ShiftReg_row_10_2$1_0/gc[9] ShiftReg_row_10_2$1_0/gc[10] d_out ShiftReg_row_10_2$1_0/PHI_1
+ ShiftReg_row_10_2$1_0/PHI_2 ShiftReg_row_10_2$1_0/D_in ShiftReg_row_10_2$1_0/Q[4]
+ ShiftReg_row_10_2$1_0/Q[9] ShiftReg_row_10_2$1_0/Q[3] ShiftReg_row_10_2$1_0/Q[8]
+ ShiftReg_row_10_2$1_0/Q[5] ShiftReg_row_10_2$1_0/Q[7] ShiftReg_row_10_2$1_0/Q[6]
+ ShiftReg_row_10_2$1_0/Q[1] ShiftReg_row_10_2$1_0/Q[2] ShiftReg_row_10_2$1_0/EN VSUBS
+ ShiftReg_row_10_2$1
Xswmatrix_Tgate_0 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[7] BUS[7]
+ swmatrix_Tgate
Xswmatrix_Tgate_1 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[9] BUS[9]
+ swmatrix_Tgate
Xswmatrix_Tgate_2 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[10] BUS[10]
+ swmatrix_Tgate
Xswmatrix_Tgate_3 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[8] BUS[8]
+ swmatrix_Tgate
Xswmatrix_Tgate_4 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[3] BUS[3]
+ swmatrix_Tgate
Xswmatrix_Tgate_5 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[5] BUS[5]
+ swmatrix_Tgate
Xswmatrix_Tgate_6 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[6] BUS[6]
+ swmatrix_Tgate
Xswmatrix_Tgate_7 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[4] BUS[4]
+ swmatrix_Tgate
Xswmatrix_Tgate_8 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[2] BUS[2]
+ swmatrix_Tgate
Xswmatrix_Tgate_9 VSUBS swmatrix_Tgate_9/VDD pin ShiftReg_row_10_2$1_0/gc[1] BUS[1]
+ swmatrix_Tgate
.ends

