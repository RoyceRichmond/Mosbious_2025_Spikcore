magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l34d0 >>
<< l21d0 >>
<< labels >>
rlabel l34d10 -0.0445 -0.178 -0.0445 -0.178 0 out
rlabel l34d10 0.017 -0.175 0.017 -0.175 0 in
rlabel l34d10 0.0305 -0.4175 0.0305 -0.4175 0 vss
rlabel l34d10 0.018 0.11 0.018 0.11 0 vdd
use pfetx241 pfetx241_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx243 nfetx243_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx243 via_devx243_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
<< end >>
