** sch_path: /foss/designs/Mosbious_2025_spiking4all/designs/libs/core_TG_bootstrapped/TG_bootstrapped.sch
.subckt TG_bootstrapped vdd vss clk nclk vin vout
*.PININFO vdd:B vss:B clk:B vin:B vout:B nclk:B
M1 net3 nclk vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M2 net1 clk vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XC2 net1 net3 cap_mim_2f0fF c_width=1e-6 c_length=1e-6 m=10
M3 net2 clk net1 vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M4 net2 nclk net1 vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M5 net2 nclk vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M6 net2 clk vss vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M7 net3 clk vin vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M8 net3 nclk vin vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M9 net5 clk vss vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M10 net4 nclk vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
XC1 net4 net5 cap_mim_2f0fF c_width=1e-6 c_length=1e-6 m=10
M11 net6 clk net5 vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M12 net6 nclk net5 vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M13 net6 nclk vdd vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M14 net6 clk vdd vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M15 vin clk net4 vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M16 vin nclk net4 vdd pfet_03v3 L=0.28u W=0.42u nf=1 m=1
M17 vout net2 vin vss nfet_03v3 L=0.28u W=0.42u nf=1 m=1
M18 vout net6 vin vdd pfet_03v3 L=0.28u W=0.84u nf=1 m=1
.ends
