* NGSPICE file created from DFF_10_row.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt DFF_2phase_1$1 gated_control PHI_1 D EN PHI_2 VDD Q VSS
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q PHI_2 Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1_0 EN Q VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1_0/I
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0/I VDD VSS gated_control
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends

.subckt DFF_10_row VDD VSS PHI_1 PHI_2 D_in Q[10] Q[4] Q[9] Q[3] Q[8] Q[5] Q[7] Q[6]
+ Q[1] Q[2] EN
XDFF_2phase_1$1_0 DFF_2phase_1$1_0/gated_control PHI_1 Q[9] EN PHI_2 DFF_2phase_1$1_9/VDD
+ DFF_2phase_1$1_0/Q VSS DFF_2phase_1$1
XDFF_2phase_1$1_1 DFF_2phase_1$1_1/gated_control PHI_1 Q[8] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[9] VSS DFF_2phase_1$1
XDFF_2phase_1$1_2 DFF_2phase_1$1_2/gated_control PHI_1 Q[7] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[8] VSS DFF_2phase_1$1
XDFF_2phase_1$1_3 DFF_2phase_1$1_3/gated_control PHI_1 Q[6] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[7] VSS DFF_2phase_1$1
XDFF_2phase_1$1_4 DFF_2phase_1$1_4/gated_control PHI_1 Q[5] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[6] VSS DFF_2phase_1$1
XDFF_2phase_1$1_5 DFF_2phase_1$1_5/gated_control PHI_1 Q[4] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[5] VSS DFF_2phase_1$1
XDFF_2phase_1$1_6 DFF_2phase_1$1_6/gated_control PHI_1 Q[3] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[4] VSS DFF_2phase_1$1
XDFF_2phase_1$1_7 DFF_2phase_1$1_7/gated_control PHI_1 Q[2] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[3] VSS DFF_2phase_1$1
XDFF_2phase_1$1_8 DFF_2phase_1$1_8/gated_control PHI_1 D_in EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[1] VSS DFF_2phase_1$1
XDFF_2phase_1$1_9 DFF_2phase_1$1_9/gated_control PHI_1 Q[1] EN PHI_2 DFF_2phase_1$1_9/VDD
+ Q[2] VSS DFF_2phase_1$1
.ends

