magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l34d0 >>
<< l36d0 >>
<< l38d0 >>
<< l42d0 >>
<< l35d0 >>
<< end >>
