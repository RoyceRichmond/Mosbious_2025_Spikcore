* Extracted by KLayout with GF180MCU LVS runset on : 27/08/2025 16:44

.SUBCKT not
M$1 vdd out in vdd pfet_03v3 L=0.35U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$2 vss out in vss nfet_03v3 L=0.28U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS not
