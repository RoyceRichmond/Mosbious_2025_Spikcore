magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l34d0 >>
<< l21d0 >>
<< l36d0 >>
<< l32d0 >>
<< labels >>
rlabel l34d10 -0.2375 -0.177 -0.2375 -0.177 0 out
rlabel l34d10 0.0135 -0.179 0.0135 -0.179 0 cntrl
rlabel l34d10 -0.1155 -0.1735 -0.1155 -0.1735 0 in
rlabel l34d10 -0.0945 0.108 -0.0945 0.108 0 vdd
rlabel l34d10 -0.0855 -0.4165 -0.0855 -0.4165 0 vss
use via_devx2428 via_devx2428_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2428 via_devx2428_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2428 via_devx2428_3
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2428 via_devx2428_4
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2418 nfetx2418_1
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use pfetx2413 pfetx2413_1
timestamp 1757365861
transform -1 0 0 0 1 0
box 0 0 0 0
use via_devx2429 via_devx2429_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx2429 via_devx2429_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx2418 nfetx2418_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use pfetx2413 pfetx2413_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
<< end >>
