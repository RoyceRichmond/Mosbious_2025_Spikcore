magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
rect -1 -1 0 1
<< l34d0 >>
rect -1 -1 0 0
<< l22d0 >>
<< l31d0 >>
<< l21d0 >>
<< l36d0 >>
<< l42d0 >>
<< l32d0 >>
<< labels >>
rlabel l34d10 -0.4545 0.6695 -0.4545 0.6695 0 vdd
rlabel l34d10 -0.192 -0.24 -0.192 -0.24 0 vp
rlabel l34d10 0.1765 -0.2385 0.1765 -0.2385 0 vn
rlabel l34d10 -0.2815 -0.4215 -0.2815 -0.4215 0 vss
rlabel l42d10 0.24 0.257 0.24 0.257 0 vout
use nfetx246 nfetx246_1
timestamp 1757365861
transform 0 -1 -1 1 0 0
box 0 0 1 0
use via_devx246 via_devx246_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx247 via_devx247_1
timestamp 1757365861
transform 1 0 0 0 1 1
box 0 0 0 0
use via_devx247 via_devx247_2
timestamp 1757365861
transform 1 0 0 0 1 1
box 0 0 0 0
use via_devx246 via_devx246_3
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_4
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx247 nfetx247_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx247 nfetx247_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx247 via_devx247_3
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use nfetx248 nfetx248_1
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_5
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx247 via_devx247_4
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_6
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use nfetx248 nfetx248_2
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_7
timestamp 1757365861
transform 0 -1 -1 1 0 0
box 0 0 0 0
use via_devx246 via_devx246_8
timestamp 1757365861
transform 1 0 -1 0 1 1
box 0 0 0 0
use via_devx247 via_devx247_5
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx248 via_devx248_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use via_devx246 via_devx246_9
timestamp 1757365861
transform 1 0 -1 0 1 0
box 0 0 0 0
use via_devx247 via_devx247_6
timestamp 1757365861
transform 0 -1 -1 1 0 0
box 0 0 0 0
use pfetx245 pfetx245_1
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
use pfetx245 pfetx245_2
timestamp 1757365861
transform 1 0 0 0 1 0
box 0 0 0 0
<< end >>
