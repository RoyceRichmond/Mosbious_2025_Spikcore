magic
tech gf180mcu
timestamp 1757365861
<< checkpaint >>
<< l42d0 >>
<< l40d0 >>
<< l46d0 >>
<< end >>
