* NGSPICE file created from top.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$5 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1$3 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt NO_ClkGen$1 clk phi_2 phi_1 vdd vss
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_11 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_11/I vdd vss
+ phi_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_12 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_12/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$5_13/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_13 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_13/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$5_13/ZN vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_14 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_14/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$5_12/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_15 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_9/ZN vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$5_14/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_0/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_1/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_17 clk vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_16/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_16 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_16/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$5_16/ZN vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_1 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_1/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_7/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_2 phi_2 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_0/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_3 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_3/I vdd vss phi_2
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_5 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_5/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_5/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_4 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_4/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_5/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_6 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_6/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_4/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_7 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_7/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_6/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_8 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_8/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_9/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_9 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_9/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_9/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$3_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_13/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$5_16/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_3/I vdd vss gf180mcu_fd_sc_mcu9t5v0__nand2_1$3
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$3_1 gf180mcu_fd_sc_mcu9t5v0__inv_1$5_5/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$5_16/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_11/I vdd vss gf180mcu_fd_sc_mcu9t5v0__nand2_1$3
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$5_10 phi_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5_8/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$5
.ends

.subckt nfet$36 a_1158_0# a_n84_n2# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_1158_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=5.6u
.ends

.subckt nfet$34 a_n84_n2# a_374_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_374_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=1.68u
.ends

.subckt pfet$19 a_150_0# a_38_n60# a_n92_0# w_n230_n138#
X0 a_150_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.286p pd=2.18u as=0.286p ps=2.18u w=0.44u l=0.56u
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=6u c_length=5u
.ends

.subckt pfet$20 a_38_n60# a_n92_0# a_318_0# w_n230_n138#
X0 a_318_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=1.4u
.ends

.subckt nfet$35 a_n84_n2# a_194_0# dw_n710_n726# a_38_n132# w_n710_n726#
X0 a_194_0# a_38_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.78u
.ends

.subckt nfet$33 a_150_0# dw_n710_n726# a_n84_0# a_38_n132# w_n710_n726#
X0 a_150_0# a_38_n132# a_n84_0# w_n710_n726# nfet_03v3 ad=0.2684p pd=2.1u as=0.2684p ps=2.1u w=0.44u l=0.56u
.ends

.subckt AH_neuron$1 vdd Current_in v_bias vout vss
Xnfet$36_0 m1_335_n170# Current_in nfet$36_0/dw_n710_n726# v_bias vss nfet$36
Xnfet$34_0 m1_335_n170# vss nfet$36_0/dw_n710_n726# vout vss nfet$34
Xpfet$19_0 vdd Current_in m2_381_1901# vdd pfet$19
Xcap_mim$3_0 Current_in vout cap_mim$3
Xpfet$20_0 m2_381_1901# vout vdd vdd pfet$20
Xnfet$35_0 vout vss nfet$36_0/dw_n710_n726# m2_381_1901# vss nfet$35
Xnfet$33_0 vss nfet$36_0/dw_n710_n726# m2_381_1901# Current_in vss nfet$33
.ends

.subckt nfet$47 a_280_0# a_158_0# a_38_n60# a_n84_0#
X0 a_158_0# a_38_n60# a_n84_0# a_280_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.6u
.ends

.subckt nfet$45 a_216_0# a_30_280# a_n84_0# a_94_0#
X0 a_94_0# a_30_280# a_n84_0# a_216_0# nfet_03v3 ad=0.671p pd=3.42u as=0.671p ps=3.42u w=1.1u l=0.28u
.ends

.subckt nfet$43 a_216_0# a_n84_0# a_94_0# a_30_480#
X0 a_94_0# a_30_480# a_n84_0# a_216_0# nfet_03v3 ad=1.281p pd=5.42u as=1.281p ps=5.42u w=2.1u l=0.28u
.ends

.subckt nfet$41 a_216_0# a_30_560# a_n84_0# a_94_0#
X0 a_94_0# a_30_560# a_n84_0# a_216_0# nfet_03v3 ad=1.525p pd=6.22u as=1.525p ps=6.22u w=2.5u l=0.28u
.ends

.subckt pfet$28 a_n92_0# a_94_0# a_28_220# w_n230_n138#
X0 a_94_0# a_28_220# a_n92_0# w_n230_n138# pfet_03v3 ad=0.52p pd=2.9u as=0.52p ps=2.9u w=0.8u l=0.28u
.ends

.subckt pfet$26 a_n92_0# a_94_0# a_28_260# w_n230_n138#
X0 a_94_0# a_28_260# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$48 a_n84_n2# a_560_n2# a_38_n60# a_438_0#
X0 a_438_0# a_38_n60# a_n84_n2# a_560_n2# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=2u
.ends

.subckt nfet$46 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$44 a_32_260# a_98_0# a_n84_0# a_220_0#
X0 a_98_0# a_32_260# a_n84_0# a_220_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
.ends

.subckt pfet$29 a_38_n60# a_n92_0# a_198_0# w_n230_n138#
X0 a_198_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.5u as=1.04p ps=4.5u w=1.6u l=0.8u
.ends

.subckt nfet$42 a_216_0# a_n84_0# a_94_0# a_30_460#
X0 a_94_0# a_30_460# a_n84_0# a_216_0# nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$27 a_238_0# a_38_n60# a_n92_0# w_n230_n138#
X0 a_238_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=1u
.ends

.subckt pfet$25 a_28_144# w_n232_n142# a_94_0# a_n92_n2#
X0 a_94_0# a_28_144# a_n92_n2# w_n232_n142# pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
.ends

.subckt schmitt_trigger vdd out in vss
Xnfet$47_0 vss vss vdd m3_n9961_n6054# nfet$47
Xnfet$45_0 vss m3_n8390_n6986# m2_n8799_n7122# vdd nfet$45
Xnfet$43_0 vss m2_n8799_n7122# vss in nfet$43
Xnfet$41_0 vss in m3_n9961_n6054# m3_n8390_n6986# nfet$41
Xpfet$28_0 m2_n8799_n7122# vdd m2_n8799_n7122# vdd pfet$28
Xpfet$26_0 m3_n9961_n6054# vdd vss vdd pfet$26
Xpfet$26_1 out vdd m3_n9961_n6054# vdd pfet$26
Xnfet$48_0 m3_n8390_n6986# vss vdd vss nfet$48
Xnfet$46_0 vss m3_n9961_n6054# out vss nfet$46
Xnfet$44_0 m3_n9961_n6054# vdd m3_n8390_n6986# vss nfet$44
Xpfet$29_0 vss m3_n8390_n6986# vdd vdd pfet$29
Xnfet$42_0 vss m2_n8799_n7122# m3_n8390_n6986# in nfet$42
Xpfet$27_0 vdd out m3_n9961_n6054# vdd pfet$27
Xpfet$25_0 in vdd vdd m3_n9961_n6054# pfet$25
.ends

.subckt cap_mim$2$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
.ends

.subckt nfet$33$1 a_216_0# a_30_172# a_n84_0# a_94_0#
X0 a_94_0# a_30_172# a_n84_0# a_216_0# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt pfet$19$1 a_38_n60# a_n92_0# a_206_0# w_n230_n138#
X0 a_206_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
.ends

.subckt nfet$32$1 a_328_0# a_38_n60# a_n84_0# a_206_0#
X0 a_206_0# a_38_n60# a_n84_0# a_328_0# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
.ends

.subckt pfet$21$1 a_2190_0# a_1250_0# a_1062_0# a_3130_0# a_3694_0# a_2942_0# a_2002_0#
+ a_2754_0# a_2566_0# a_2378_0# a_1814_0# a_1626_0# a_1438_0# a_602_n60# a_414_n60#
+ a_226_n60# a_2670_n60# a_3506_0# a_3318_0# a_2482_n60# a_2294_n60# a_3610_n60# a_3422_n60#
+ a_3234_n60# a_2858_n60# a_38_n60# a_3046_n60# a_n92_0# a_310_0# a_122_0# a_874_0#
+ a_686_0# a_498_0# a_1730_n60# a_1542_n60# a_790_n60# a_1918_n60# a_1354_n60# a_1166_n60#
+ a_2106_n60# a_978_n60# w_n230_n138#
X0 a_2378_0# a_2294_n60# a_2190_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X1 a_2942_0# a_2858_n60# a_2754_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X2 a_3694_0# a_3610_n60# a_3506_0# w_n230_n138# pfet_03v3 ad=2.028p pd=7.54u as=0.8112p ps=3.64u w=3.12u l=0.42u
X3 a_2566_0# a_2482_n60# a_2378_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X4 a_2754_0# a_2670_n60# a_2566_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X5 a_310_0# a_226_n60# a_122_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X6 a_498_0# a_414_n60# a_310_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X7 a_686_0# a_602_n60# a_498_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X8 a_2190_0# a_2106_n60# a_2002_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X9 a_2002_0# a_1918_n60# a_1814_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X10 a_1250_0# a_1166_n60# a_1062_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X11 a_1438_0# a_1354_n60# a_1250_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X12 a_1626_0# a_1542_n60# a_1438_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X13 a_1814_0# a_1730_n60# a_1626_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X14 a_122_0# a_38_n60# a_n92_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=2.028p ps=7.54u w=3.12u l=0.42u
X15 a_1062_0# a_978_n60# a_874_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X16 a_874_0# a_790_n60# a_686_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X17 a_3130_0# a_3046_n60# a_2942_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X18 a_3318_0# a_3234_n60# a_3130_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X19 a_3506_0# a_3422_n60# a_3318_0# w_n230_n138# pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
.ends

.subckt pfet$18$1 a_n92_0# a_38_n136# a_206_0# w_n230_n138#
X0 a_206_0# a_38_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
.ends

.subckt nfet$31$1 a_328_0# a_n84_0# a_38_n132# a_206_0#
X0 a_206_0# a_38_n132# a_n84_0# a_328_0# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
.ends

.subckt nfet$34$1 a_2190_0# a_414_n132# a_1250_0# a_1062_0# a_2670_n132# a_790_n132#
+ a_1542_n132# a_2942_0# a_2002_0# a_2754_0# a_2566_0# a_2378_0# a_1814_0# a_1626_0#
+ a_2858_n132# a_1438_0# a_2106_n132# a_978_n132# a_226_n132# a_3064_0# a_2482_n132#
+ a_310_0# a_122_0# a_n84_0# a_1354_n132# a_602_n132# a_874_0# a_686_0# a_498_0# a_38_n132#
+ a_1730_n132# a_2294_n132# a_1918_n132# a_1166_n132#
X0 a_2378_0# a_2294_n132# a_2190_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X1 a_2566_0# a_2482_n132# a_2378_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X2 a_2754_0# a_2670_n132# a_2566_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X3 a_310_0# a_226_n132# a_122_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X4 a_498_0# a_414_n132# a_310_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X5 a_686_0# a_602_n132# a_498_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X6 a_2190_0# a_2106_n132# a_2002_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X7 a_2002_0# a_1918_n132# a_1814_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X8 a_1250_0# a_1166_n132# a_1062_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X9 a_1438_0# a_1354_n132# a_1250_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X10 a_1626_0# a_1542_n132# a_1438_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X11 a_1814_0# a_1730_n132# a_1626_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X12 a_122_0# a_38_n132# a_n84_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=2.38815p ps=9.05u w=3.915u l=0.42u
X13 a_1062_0# a_978_n132# a_874_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X14 a_874_0# a_790_n132# a_686_0# a_3064_0# nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X15 a_2942_0# a_2858_n132# a_2754_0# a_3064_0# nfet_03v3 ad=2.38815p pd=9.05u as=1.0179p ps=4.435u w=3.915u l=0.42u
.ends

.subckt pfet$20$1 a_28_284# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_284# a_n92_0# w_n230_n138# pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
.ends

.subckt TG_bootstrapped clk vss vin nclk vout vdd
Xcap_mim$2$1_0 m4_6353_n3083# m5_6577_n2963# cap_mim$2$1
Xcap_mim$2$1_1 m4_6354_2903# m5_6578_3023# cap_mim$2$1
Xnfet$33$1_0 vss nclk m5_6577_n2963# vss nfet$33$1
Xnfet$33$1_1 vss clk m4_6354_2903# vss nfet$33$1
Xpfet$19$1_0 nclk m5_6577_n2963# vin vdd pfet$19$1
Xnfet$32$1_0 vss clk m5_6577_n2963# vin nfet$32$1
Xpfet$19$1_1 clk vss m1_5676_n176# vdd pfet$19$1
Xnfet$32$1_1 vss clk m4_6353_n3083# m1_5676_n176# nfet$32$1
Xpfet$19$1_2 nclk m5_6578_3023# vin vdd pfet$19$1
Xnfet$32$1_2 vss clk m5_6578_3023# vin nfet$32$1
Xpfet$19$1_3 clk vdd m3_6686_2072# vdd pfet$19$1
Xnfet$32$1_3 vss clk m4_6354_2903# m3_6686_2072# nfet$32$1
Xpfet$21$1_0 vout vin vout vin vout vout vin vin vout vin vout vin vout m3_6686_2072#
+ m3_6686_2072# m3_6686_2072# m3_6686_2072# vin vout m3_6686_2072# m3_6686_2072# m3_6686_2072#
+ m3_6686_2072# m3_6686_2072# m3_6686_2072# m3_6686_2072# m3_6686_2072# vout vout
+ vin vin vout vin m3_6686_2072# m3_6686_2072# m3_6686_2072# m3_6686_2072# m3_6686_2072#
+ m3_6686_2072# m3_6686_2072# m3_6686_2072# vdd pfet$21$1
Xpfet$18$1_0 m4_6353_n3083# nclk m1_5676_n176# vdd pfet$18$1
Xnfet$31$1_0 vss vss nclk m1_5676_n176# nfet$31$1
Xpfet$18$1_1 m4_6354_2903# nclk m3_6686_2072# vdd pfet$18$1
Xnfet$31$1_1 vss vdd nclk m3_6686_2072# nfet$31$1
Xnfet$34$1_0 vout m1_5676_n176# vin vout m1_5676_n176# m1_5676_n176# m1_5676_n176#
+ vout vin vin vout vin vout vin m1_5676_n176# vout m1_5676_n176# m1_5676_n176# m1_5676_n176#
+ vss m1_5676_n176# vout vin vout m1_5676_n176# m1_5676_n176# vin vout vin m1_5676_n176#
+ m1_5676_n176# m1_5676_n176# m1_5676_n176# m1_5676_n176# nfet$34$1
Xpfet$20$1_0 clk m4_6353_n3083# vdd vdd pfet$20$1
Xpfet$20$1_1 nclk m5_6578_3023# vdd vdd pfet$20$1
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$7 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$1 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt En_clk_din clk d_in data_in clock vdd vss Enable
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$7_0 Enable vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$7_0/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$7
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$7_1 Enable vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$7_1/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$7
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$7_0/ZN d_in vdd
+ vss data_in vdd vss gf180mcu_fd_sc_mcu9t5v0__and2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_1 gf180mcu_fd_sc_mcu9t5v0__inv_1$7_1/ZN clk vdd
+ vss clock vdd vss gf180mcu_fd_sc_mcu9t5v0__and2_1$1
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1$4 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$8 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt NO_ClkGen clk phi_2 phi_1 vdd vss
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$4_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_13/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$8_16/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_3/I vdd vss gf180mcu_fd_sc_mcu9t5v0__nand2_1$4
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_10 phi_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_8/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$4_1 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_5/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$8_16/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_11/I vdd vss gf180mcu_fd_sc_mcu9t5v0__nand2_1$4
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_11 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_11/I vdd vss
+ phi_1 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_13 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_13/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$8_13/ZN vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_12 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_12/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$8_13/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_14 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_14/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$8_12/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_15 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_9/ZN vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$8_14/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_16 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_16/I vdd vss
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$8_16/ZN vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_17 clk vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_16/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_0/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_1/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_2 phi_2 vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_0/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_1 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_1/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_7/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_3 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_3/I vdd vss phi_2
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_4 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_4/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_5/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_5 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_5/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_5/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_6 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_6/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_4/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_7 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_7/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_6/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_8 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_8/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_9/I
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$8_9 gf180mcu_fd_sc_mcu9t5v0__inv_1$8_9/I vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8_9/ZN
+ vdd vss gf180mcu_fd_sc_mcu9t5v0__inv_1$8
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$10 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt pfet$18 a_1534_0# a_2174_0# a_1054_0# a_734_0# a_828_n136# a_28_n136# a_2588_n136#
+ a_1694_0# a_254_0# a_1628_n136# a_894_0# a_188_n136# a_988_n136# a_2814_0# a_2748_n136#
+ a_1788_n136# a_2334_0# a_348_n136# a_1214_0# a_1148_n136# a_1854_0# a_414_0# a_2108_n136#
+ a_2494_0# a_n92_0# a_1948_n136# a_1374_0# a_94_0# a_574_0# a_508_n136# a_2268_n136#
+ a_1308_n136# a_2014_0# a_668_n136# a_2428_n136# a_1468_n136# a_2654_0# w_n230_n138#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1 a_2654_0# a_2588_n136# a_2494_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X2 a_734_0# a_668_n136# a_574_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X3 a_2494_0# a_2428_n136# a_2334_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X4 a_254_0# a_188_n136# a_94_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X5 a_574_0# a_508_n136# a_414_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X6 a_2014_0# a_1948_n136# a_1854_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X7 a_1534_0# a_1468_n136# a_1374_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X8 a_1374_0# a_1308_n136# a_1214_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X9 a_1054_0# a_988_n136# a_894_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X10 a_2814_0# a_2748_n136# a_2654_0# w_n230_n138# pfet_03v3 ad=2.6p pd=9.3u as=1.04p ps=4.52u w=4u l=0.28u
X11 a_894_0# a_828_n136# a_734_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X12 a_2334_0# a_2268_n136# a_2174_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X13 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=2.6p ps=9.3u w=4u l=0.28u
X14 a_2174_0# a_2108_n136# a_2014_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X15 a_414_0# a_348_n136# a_254_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X16 a_1854_0# a_1788_n136# a_1694_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X17 a_1694_0# a_1628_n136# a_1534_0# w_n230_n138# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
.ends

.subckt nfet$31 vss a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_830_n132#
+ a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_350_n132#
X0 a_734_0# a_670_n132# a_574_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X3 a_894_0# a_830_n132# a_734_0# vss nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.28u
X4 a_94_0# a_30_n132# a_n84_0# vss nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.28u
X5 a_414_0# a_350_n132# a_254_0# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
.ends

.subckt swmatrix_Tgate$1 VSS VDD T1 gated_control T2
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$10_0 gated_control VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$10
Xpfet$18_0 T1 T1 T2 T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN T2 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ T1 T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN T1 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ T2 T2 T1 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN T2 gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN
+ gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN gf180mcu_fd_sc_mcu9t5v0__inv_1$10_0/ZN T2
+ VDD pfet$18
Xnfet$31_0 VSS T2 gated_control T1 T1 gated_control gated_control T2 gated_control
+ T1 T2 gated_control T1 gated_control nfet$31
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1$5 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$2 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$9 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt DFF_2phase_1$2 gated_control PHI_1 D PHI_2 EN Q VDD VSS
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$5_0 EN Q VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$9_0/I
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1$5
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$2_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$2_1/Q PHI_2 Q
+ VDD VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1$2
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$2_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$2_1/Q
+ VDD VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1$2
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$9_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$9_0/I VDD VSS gated_control
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$9
.ends

.subckt ShiftReg_row_10_2$1 gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8] gc[9]
+ gc[10] Q[10] PHI_1 PHI_2 Q[4] Q[9] Q[3] Q[8] Q[5] Q[7] Q[6] Q[1] Q[2] EN D_in VSS
+ VDD
XDFF_2phase_1$2_8 gc[1] PHI_1 D_in PHI_2 EN Q[1] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_9 gc[2] PHI_1 Q[1] PHI_2 EN Q[2] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_0 gc[10] PHI_1 Q[9] PHI_2 EN Q[10] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_1 gc[9] PHI_1 Q[8] PHI_2 EN Q[9] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_2 gc[8] PHI_1 Q[7] PHI_2 EN Q[8] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_3 gc[7] PHI_1 Q[6] PHI_2 EN Q[7] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_4 gc[6] PHI_1 Q[5] PHI_2 EN Q[6] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_5 gc[5] PHI_1 Q[4] PHI_2 EN Q[5] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_6 gc[4] PHI_1 Q[3] PHI_2 EN Q[4] VDD VSS DFF_2phase_1$2
XDFF_2phase_1$2_7 gc[3] PHI_1 Q[2] PHI_2 EN Q[3] VDD VSS DFF_2phase_1$2
.ends

.subckt swmatrix_row_10 pin BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] d_out ShiftReg_row_10_2$1_0/EN ShiftReg_row_10_2$1_0/D_in ShiftReg_row_10_2$1_0/PHI_2
+ VSUBS ShiftReg_row_10_2$1_0/PHI_1 swmatrix_Tgate$1_9/VDD
Xswmatrix_Tgate$1_0 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[7] BUS[7]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_1 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[9] BUS[9]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_2 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[10]
+ BUS[10] swmatrix_Tgate$1
Xswmatrix_Tgate$1_3 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[8] BUS[8]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_4 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[3] BUS[3]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_5 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[5] BUS[5]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_6 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[6] BUS[6]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_7 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[4] BUS[4]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_8 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[2] BUS[2]
+ swmatrix_Tgate$1
Xswmatrix_Tgate$1_9 VSUBS swmatrix_Tgate$1_9/VDD pin ShiftReg_row_10_2$1_0/gc[1] BUS[1]
+ swmatrix_Tgate$1
XShiftReg_row_10_2$1_0 ShiftReg_row_10_2$1_0/gc[1] ShiftReg_row_10_2$1_0/gc[2] ShiftReg_row_10_2$1_0/gc[3]
+ ShiftReg_row_10_2$1_0/gc[4] ShiftReg_row_10_2$1_0/gc[5] ShiftReg_row_10_2$1_0/gc[6]
+ ShiftReg_row_10_2$1_0/gc[7] ShiftReg_row_10_2$1_0/gc[8] ShiftReg_row_10_2$1_0/gc[9]
+ ShiftReg_row_10_2$1_0/gc[10] d_out ShiftReg_row_10_2$1_0/PHI_1 ShiftReg_row_10_2$1_0/PHI_2
+ ShiftReg_row_10_2$1_0/Q[4] ShiftReg_row_10_2$1_0/Q[9] ShiftReg_row_10_2$1_0/Q[3]
+ ShiftReg_row_10_2$1_0/Q[8] ShiftReg_row_10_2$1_0/Q[5] ShiftReg_row_10_2$1_0/Q[7]
+ ShiftReg_row_10_2$1_0/Q[6] ShiftReg_row_10_2$1_0/Q[1] ShiftReg_row_10_2$1_0/Q[2]
+ ShiftReg_row_10_2$1_0/EN ShiftReg_row_10_2$1_0/D_in VSUBS swmatrix_Tgate$1_9/VDD
+ ShiftReg_row_10_2$1
.ends

.subckt swmatrix_24_by_10 PIN[1] PIN[2] PIN[3] PIN[4] PIN[5] PIN[6] PIN[7] PIN[8]
+ PIN[9] PIN[10] PIN[11] PIN[12] PIN[13] PIN[14] PIN[15] PIN[16] PIN[17] PIN[21] PIN[18]
+ PIN[19] PIN[20] PIN[22] PIN[23] PIN[24] D_out clk d_in BUS[1] BUS[2] BUS[3] BUS[4]
+ BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] swmatrix_row_10_0[6]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[20]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[12]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[1]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[18]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[21]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[13]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[2]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[8]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[22]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[14]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[3]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[15]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[4]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[10]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[7]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[16]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[5]/swmatrix_Tgate$1_9/VDD swmatrix_row_10_0[9]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[11]/swmatrix_Tgate$1_9/VDD vdd Enable NO_ClkGen_0/phi_2 swmatrix_row_10_0[0]/ShiftReg_row_10_2$1_0/PHI_1
+ swmatrix_row_10_0[0]/swmatrix_Tgate$1_9/VDD vss swmatrix_row_10_0[17]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10_0[19]/swmatrix_Tgate$1_9/VDD
XEn_clk_din_0 clk d_in En_clk_din_0/data_in NO_ClkGen_0/clk vdd vss Enable En_clk_din
XNO_ClkGen_0 NO_ClkGen_0/clk NO_ClkGen_0/phi_2 NO_ClkGen_0/phi_1 vdd vss NO_ClkGen
Xswmatrix_row_10_0[0] PIN[24] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] D_out Enable swmatrix_row_10_0[0]/ShiftReg_row_10_2$1_0/D_in NO_ClkGen_0/phi_2
+ vss swmatrix_row_10_0[0]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[0]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[1] PIN[23] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[1]/d_out Enable swmatrix_row_10_0[1]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[1]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[1]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[2] PIN[22] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[2]/d_out Enable swmatrix_row_10_0[2]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[2]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[2]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[3] PIN[21] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[3]/d_out Enable swmatrix_row_10_0[3]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[3]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[3]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[4] PIN[20] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[4]/d_out Enable swmatrix_row_10_0[4]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[4]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[4]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[5] PIN[19] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[5]/d_out Enable swmatrix_row_10_0[5]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[5]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[5]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[6] PIN[18] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[6]/d_out Enable swmatrix_row_10_0[6]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[6]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[6]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[7] PIN[17] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[7]/d_out Enable swmatrix_row_10_0[7]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[7]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[7]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[8] PIN[16] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[8]/d_out Enable swmatrix_row_10_0[8]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[8]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[8]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[9] PIN[15] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[9]/d_out Enable swmatrix_row_10_0[9]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[9]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[9]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[10] PIN[14] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[10]/d_out Enable swmatrix_row_10_0[10]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[10]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[10]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[11] PIN[13] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[11]/d_out Enable swmatrix_row_10_0[11]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[11]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[11]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[12] PIN[12] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[12]/d_out Enable swmatrix_row_10_0[12]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[12]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[12]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[13] PIN[11] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[13]/d_out Enable swmatrix_row_10_0[13]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[13]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[13]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[14] PIN[10] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[14]/d_out Enable swmatrix_row_10_0[14]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[14]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[14]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[15] PIN[9] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[15]/d_out Enable swmatrix_row_10_0[15]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[15]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[15]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[16] PIN[8] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[16]/d_out Enable swmatrix_row_10_0[16]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[16]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[16]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[17] PIN[7] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[17]/d_out Enable swmatrix_row_10_0[17]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[17]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[17]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[18] PIN[6] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[18]/d_out Enable swmatrix_row_10_0[18]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[18]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[18]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[19] PIN[5] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[19]/d_out Enable swmatrix_row_10_0[19]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[19]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[19]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[20] PIN[4] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[20]/d_out Enable swmatrix_row_10_0[20]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[20]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[20]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[21] PIN[3] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[21]/d_out Enable swmatrix_row_10_0[21]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[21]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[21]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[22] PIN[2] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[22]/d_out Enable swmatrix_row_10_0[22]/ShiftReg_row_10_2$1_0/D_in
+ NO_ClkGen_0/phi_2 vss swmatrix_row_10_0[22]/ShiftReg_row_10_2$1_0/PHI_1 swmatrix_row_10_0[22]/swmatrix_Tgate$1_9/VDD
+ swmatrix_row_10
Xswmatrix_row_10_0[23] PIN[1] BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8]
+ BUS[9] BUS[10] swmatrix_row_10_0[23]/d_out Enable En_clk_din_0/data_in NO_ClkGen_0/phi_2
+ vss NO_ClkGen_0/phi_1 vdd swmatrix_row_10
.ends

.subckt pfet$23 a_28_144# w_n232_n142# a_94_0# a_n92_n2#
X0 a_94_0# a_28_144# a_n92_n2# w_n232_n142# pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
.ends

.subckt pfet$21 a_28_620# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_620# a_n92_0# w_n230_n138# pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
.ends

.subckt nfet$38 a_n84_n2# dw_n710_n726# a_30_n132# a_94_0# w_n710_n726#
X0 a_94_0# a_30_n132# a_n84_n2# w_n710_n726# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
.ends

.subckt pfet$24 a_28_n136# w_n232_n142# a_94_0# a_n92_n2#
X0 a_94_0# a_28_n136# a_n92_n2# w_n232_n142# pfet_03v3 ad=0.2822p pd=2.18u as=0.2822p ps=2.18u w=0.42u l=0.28u
.ends

.subckt pfet$22 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
.ends

.subckt nfet$39 dw_n710_n652# a_30_260# a_n84_0# a_94_0# w_n710_n652#
X0 a_94_0# a_30_260# a_n84_0# w_n710_n652# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nfet$37 dw_n710_n726# a_30_n132# a_n84_0# a_94_0# w_n710_n726#
X0 a_94_0# a_30_n132# a_n84_0# w_n710_n726# nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$40 a_n84_n2# dw_n710_n652# a_94_0# a_30_144# w_n710_n652#
X0 a_94_0# a_30_144# a_n84_n2# w_n710_n652# nfet_03v3 ad=0.2646p pd=2.1u as=0.2646p ps=2.1u w=0.42u l=0.28u
.ends

.subckt synapse vi v_ctrl v_in ve vdd v_out m1_344_2455# vss
Xpfet$23_1 m1_856_n14# vdd m1_44_2533# m1_344_2455# pfet$23
Xpfet$23_0 v_in vdd vdd m1_856_n14# pfet$23
Xpfet$23_2 m2_640_1617# vdd vdd m2_640_1617# pfet$23
Xpfet$21_0 v_ctrl v_out m1_1750_2493# vdd pfet$21
Xnfet$38_0 m1_1434_n778# nfet$40_0/dw_n710_n652# ve vss vss nfet$38
Xnfet$38_2 m1_344_2455# nfet$40_0/dw_n710_n652# m1_344_2455# vss vss nfet$38
Xnfet$38_1 m1_856_n14# nfet$40_0/dw_n710_n652# v_in vss vss nfet$38
Xpfet$24_0 vi vdd vdd m1_44_2533# pfet$24
Xpfet$22_0 m2_640_1617# m1_1750_2493# vdd vdd pfet$22
Xnfet$39_0 nfet$40_0/dw_n710_n652# m1_344_2455# m1_2266_n82# vss vss nfet$39
Xnfet$37_0 nfet$40_0/dw_n710_n652# v_ctrl v_out m1_2266_n82# vss nfet$37
Xnfet$40_0 m2_640_1617# nfet$40_0/dw_n710_n652# m1_1434_n778# v_in vss nfet$40
.ends

.subckt AH_neuron vdd Current_in v_bias vout vss
Xnfet$36_0 m1_335_n170# Current_in nfet$36_0/dw_n710_n726# v_bias vss nfet$36
Xnfet$34_0 m1_335_n170# vss nfet$36_0/dw_n710_n726# vout vss nfet$34
Xpfet$19_0 vdd Current_in m2_381_1901# vdd pfet$19
Xcap_mim$3_0 Current_in vout cap_mim$3
Xpfet$20_0 m2_381_1901# vout vdd vdd pfet$20
Xnfet$35_0 vout vss nfet$36_0/dw_n710_n726# m2_381_1901# vss nfet$35
Xnfet$33_0 vss nfet$36_0/dw_n710_n726# m2_381_1901# Current_in vss nfet$33
.ends

.subckt nfet$24 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$14 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt switch out cntrl vdd vss in
Xnfet$24_1 vss cntrl in out nfet$24
Xpfet$14_0 m2_n331_n296# cntrl vdd vdd pfet$14
Xpfet$14_1 in m2_n331_n296# out vdd pfet$14
Xnfet$24_0 vss cntrl m2_n331_n296# vss nfet$24
.ends

.subckt nfet$22 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet$23 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$21 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt pfet$13 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt ota_1stage vdd vp vn vss vout
Xnfet$22_0 vss vn m3_n530_n14# vout nfet$22
Xnfet$22_1 vss vp m3_n530_n14# m3_n314_178# nfet$22
Xnfet$23_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$23
Xnfet$23_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$23
Xnfet$21_0 m3_n1200_n476# vss vdd vdd nfet$21
Xpfet$13_0 vdd vdd m3_n314_178# m3_n314_178# pfet$13
Xpfet$13_1 vdd vdd vout m3_n314_178# pfet$13
.ends

.subckt cap_mim$2 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt pfet$16 w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$29 a_n256_n198# a_30_228# a_n84_0# a_94_0#
X0 a_94_0# a_30_228# a_n84_0# a_n256_n198# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$27 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt pfet$17 a_28_n136# a_n92_0# a_94_0# w_n352_n362#
X0 a_94_0# a_28_n136# a_n92_0# w_n352_n362# pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.28u
.ends

.subckt nfet$30 a_n256_n198# a_30_172# a_n84_0# a_94_0#
X0 a_94_0# a_30_172# a_n84_0# a_n256_n198# nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
.ends

.subckt cap_mim$1 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=9u c_length=9u
.ends

.subckt nfet$28 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt nfet$26 a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt ota_2stage vdd vp vn vss vout
Xpfet$16_0 vdd vdd m3_n314_178# m3_n314_178# pfet$16
Xpfet$16_1 vdd m3_210_178# vdd m3_n314_178# pfet$16
Xnfet$29_0 vss m3_n1200_n227# m3_n1200_n227# vss nfet$29
Xnfet$27_0 vss vp m3_210_178# m3_n530_n14# nfet$27
Xnfet$27_1 vss vn m3_n530_n14# m3_n314_178# nfet$27
Xpfet$17_0 m3_210_178# vdd vout vdd pfet$17
Xnfet$30_0 vss m3_n1200_n227# vss vout nfet$30
Xcap_mim$1_0 vout m3_210_178# cap_mim$1
Xnfet$28_0 vss m3_n1200_n227# vss m3_n530_n14# nfet$28
Xnfet$26_0 m3_n1200_n227# vss vdd vdd nfet$26
.ends

.subckt nfet$32 a_n256_n198# a_38_n60# a_n84_0# a_138_0#
X0 a_138_0# a_38_n60# a_n84_0# a_n256_n198# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$25 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$15 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt conmutator in1 in2 vdd out cntrl vss
Xnfet$25_0 vss m2_n850_n472# out in1 nfet$25
Xnfet$25_1 vss cntrl in2 out nfet$25
Xnfet$25_2 vss cntrl m2_n850_n472# vss nfet$25
Xpfet$15_0 out cntrl in1 vdd pfet$15
Xpfet$15_1 in2 m2_n850_n472# out vdd pfet$15
Xpfet$15_2 m2_n850_n472# cntrl vdd vdd pfet$15
.ends

.subckt nfet$9 a_n256_n272# a_n84_0# a_198_0# a_38_n132#
X0 a_198_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.8u
.ends

.subckt nfet$7 a_n84_n2# a_n256_n272# a_30_n132# a_94_0#
X0 a_94_0# a_30_n132# a_n84_n2# a_n256_n272# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=0.28u
.ends

.subckt nfet$8 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt nfet$10 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.3355p pd=2.32u as=0.3355p ps=2.32u w=0.55u l=0.28u
.ends

.subckt nvdiv vss vdd vspike_up vspike_down vres vref
Xnfet$9_0 vss vres vss vres nfet$9
Xnfet$7_0 vref vss vref vss nfet$7
Xnfet$7_1 vspike_up vss vspike_up m2_367_1540# nfet$7
Xnfet$7_2 vdd vss vdd vspike_up nfet$7
Xnfet$8_0 vss vspike_down vspike_down vres nfet$8
Xnfet$8_1 vss m2_367_1540# m2_367_1540# vspike_down nfet$8
Xnfet$10_0 vss vdd vdd vref nfet$10
.ends

.subckt pfet$8 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$13 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt not$1 out in vdd vss
Xpfet$8_0 out in vdd vdd pfet$8
Xnfet$13_0 vss in out vss nfet$13
.ends

.subckt pfet$7 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$12 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt switch$1 out cntrl in vdd vss
Xpfet$7_0 m2_n331_n296# cntrl vdd vdd pfet$7
Xpfet$7_1 in m2_n331_n296# out vdd pfet$7
Xnfet$12_0 vss cntrl m2_n331_n296# vss nfet$12
Xnfet$12_1 vss cntrl in out nfet$12
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt nfet$3 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$1 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt not out in vdd vss
Xnfet$3_0 vss in out vss nfet$3
Xpfet$1_0 out in vdd vdd pfet$1
.ends

.subckt pfet$4 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$5 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$3 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$4 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt nand A B Z vdd vss
Xpfet$4_0 B Z vdd vdd pfet$4
Xnfet$5_0 A Z nfet$5_0/a_94_0# vss nfet$5
Xpfet$3_0 A vdd vdd Z pfet$3
Xnfet$4_0 vss B nfet$5_0/a_94_0# vss nfet$4
.ends

.subckt nfet$19 a_98_0# a_n256_n272# a_n84_0# a_32_n132#
X0 a_98_0# a_32_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.3u
.ends

.subckt monostable vin vres phi_1 vneg vdd vss phi_2
Xcap_mim_0 not_1/in nand_0/Z cap_mim
Xcap_mim_1 not_3/in nand_1/Z cap_mim
Xnot_0 phi_2 not_0/in vdd vss not
Xnot_1 not_0/in not_1/in vdd vss not
Xnot_2 phi_1 vneg vdd vss not
Xnot_3 vneg not_3/in vdd vss not
Xnand_0 not_0/in phi_1 nand_0/Z vdd vss nand
Xnfet$19_0 vss vss not_1/in vres nfet$19
Xnfet$19_1 vss vss not_3/in vres nfet$19
Xnand_1 vneg vin nand_1/Z vdd vss nand
.ends

.subckt nfet$15 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$10 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nfet$14 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$11 a_28_n136# a_n92_0# a_94_0# w_n230_n138#
X0 a_94_0# a_28_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.28u
.ends

.subckt nor A B Z vdd vss
Xnfet$15_0 B vss Z vss nfet$15
Xpfet$10_0 B vdd Z pfet$10_0/a_94_0# pfet$10
Xnfet$14_0 vss A Z vss nfet$14
Xpfet$11_0 A pfet$10_0/a_94_0# vdd vdd pfet$11
.ends

.subckt pfet$6 a_n92_0# a_35_n136# a_108_0# w_n230_n138#
X0 a_108_0# a_35_n136# a_n92_0# w_n230_n138# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.35u
.ends

.subckt nfet$11 a_216_0# a_30_260# a_n84_0# a_94_0#
X0 a_94_0# a_30_260# a_n84_0# a_216_0# nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt conmutator$1 out in1 in2 vdd cntrl vss
Xpfet$6_0 out cntrl in1 vdd pfet$6
Xpfet$6_2 m2_n850_n472# cntrl vdd vdd pfet$6
Xpfet$6_1 in2 m2_n850_n472# out vdd pfet$6
Xnfet$11_0 vss m2_n850_n472# out in1 nfet$11
Xnfet$11_1 vss cntrl in2 out nfet$11
Xnfet$11_2 vss cntrl m2_n850_n472# vss nfet$11
.ends

.subckt nfet$17 a_n256_n198# a_30_3060# a_n84_0# a_94_0#
X0 a_94_0# a_30_3060# a_n84_0# a_n256_n198# nfet_03v3 ad=9.15p pd=31.22u as=9.15p ps=31.22u w=15u l=0.28u
.ends

.subckt nfet$18 a_2638_0# a_n84_n2# a_n256_n198# a_38_n60#
X0 a_2638_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=13u
.ends

.subckt nfet$16 a_n256_n272# a_n84_0# a_38_n132# a_138_0#
X0 a_138_0# a_38_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.5u
.ends

.subckt pfet w_n352_n286# a_n92_0# a_94_0# a_28_228#
X0 a_94_0# a_28_228# a_n92_0# w_n352_n286# pfet_03v3 ad=0.546p pd=2.98u as=0.546p ps=2.98u w=0.84u l=0.28u
.ends

.subckt nfet$1 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=1.8788p pd=7.38u as=1.8788p ps=7.38u w=3.08u l=0.28u
.ends

.subckt nfet a_n84_n2# a_n256_n198# a_1746_0# a_38_n60#
X0 a_1746_0# a_38_n60# a_n84_n2# a_n256_n198# nfet_03v3 ad=0.228p pd=1.98u as=0.228p ps=1.98u w=0.36u l=8.54u
.ends

.subckt nfet$2 a_n256_n272# a_30_n132# a_n84_0# a_94_0#
X0 a_94_0# a_30_n132# a_n84_0# a_n256_n272# nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.28u
.ends

.subckt ota_1stage$1 vdd vp vn vss vout
Xpfet_0 vdd vdd m3_n314_178# m3_n314_178# pfet
Xpfet_1 vdd vdd vout m3_n314_178# pfet
Xnfet$1_0 vss vn m3_n530_n14# vout nfet$1
Xnfet$1_1 vss vp m3_n530_n14# m3_n314_178# nfet$1
Xnfet_0 m3_n1200_n476# vss vdd vdd nfet
Xnfet$2_0 vss m3_n1200_n476# m3_n1200_n476# vss nfet$2
Xnfet$2_1 vss m3_n1200_n476# vss m3_n530_n14# nfet$2
.ends

.subckt refractory vneg vss vspike_down vdd vrefrac
Xnfet$17_0 vss ota_1stage$1_0/vp vss ota_1stage$1_0/vp nfet$17
Xnfet$18_0 vneg ota_1stage$1_0/vp vss vneg nfet$18
Xnfet$16_0 vss ota_1stage$1_0/vn vspike_down vspike_down nfet$16
Xnfet$16_1 vss ota_1stage$1_0/vn ota_1stage$1_0/vn vrefrac nfet$16
Xota_1stage$1_0 vdd ota_1stage$1_0/vp ota_1stage$1_0/vn vss vrefrac ota_1stage$1
.ends

.subckt phaseUpulse phi_fire vin vspike reward vres vdd vref vss
Xnvdiv_0 vss vdd vspike_up vspike_down vres vref nvdiv
Xnot$1_0 phi_fire phi_int vdd vss not$1
Xswitch$1_0 switch$1_0/out phi_1 vspike vdd vss switch$1
Xswitch$1_1 vrefrac phi_2 vspike vdd vss switch$1
Xmonostable_0 vin vres phi_1 vneg vdd vss phi_2 monostable
Xswitch$1_2 vref phi_int vspike vdd vss switch$1
Xnor_0 phi_1 phi_2 phi_int vdd vss nor
Xconmutator$1_0 switch$1_0/out vspike_up vdd vdd reward vss conmutator$1
Xrefractory_0 vneg vss vspike_down vdd vrefrac refractory
.ends

.subckt LIF_comp vin v_rew vout vdd vss
Xswitch_0 vmem phi_fire vdd vss vin switch
Xota_1stage_0 vdd ota_1stage_0/vp v_th vss phaseUpulse_0/vin ota_1stage
Xcap_mim$2_0 conmutator_2/out vin cap_mim$2
Xota_2stage_0 vdd vspike vin vss vmem ota_2stage
Xnfet$32_0 vss v_th vin vmem nfet$32
Xconmutator_0 vmem vss vdd ota_1stage_0/vp phi_fire vss conmutator
Xconmutator_1 v_ref vmem vdd vout phi_fire vss conmutator
Xconmutator_2 vmem v_ref vdd conmutator_2/out phi_fire vss conmutator
XphaseUpulse_0 phi_fire phaseUpulse_0/vin vspike v_rew v_th vdd v_ref vss phaseUpulse
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1$1 A1 A2 VDD VSS ZN VNW VPW
X0 ZN A2 VDD VNW pfet_05v0 ad=0.4277p pd=2.165u as=0.7238p ps=4.17u w=1.645u l=0.5u
X1 VDD A1 ZN VNW pfet_05v0 ad=0.7238p pd=4.17u as=0.4277p ps=2.165u w=1.645u l=0.5u
X2 ZN A1 a_245_69# VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.2112p ps=1.64u w=1.32u l=0.6u
X3 a_245_69# A2 VSS VPW nfet_05v0 ad=0.2112p pd=1.64u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$2 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt DFF_2phase_1 gated_control PHI_1 D EN PHI_2 Q VDD VSS
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q PHI_2 Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__nand2_1$1_0 EN Q VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$2_0/I
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__nand2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$2_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$2_0/I VDD VSS gated_control
+ VDD VSS gf180mcu_fd_sc_mcu9t5v0__inv_1$2
.ends

.subckt ShiftReg_row_10_2$2 gc[1] gc[2] gc[3] gc[4] gc[5] gc[6] gc[7] gc[8] gc[9]
+ gc[10] Q[10] PHI_2 Q[4] Q[9] Q[3] Q[8] Q[5] Q[7] Q[6] Q[1] Q[2] EN D_in PHI_1 VDD
+ VSS
XDFF_2phase_1_0 gc[10] PHI_1 Q[9] EN PHI_2 Q[10] VDD VSS DFF_2phase_1
XDFF_2phase_1_1 gc[9] PHI_1 Q[8] EN PHI_2 Q[9] VDD VSS DFF_2phase_1
XDFF_2phase_1_2 gc[8] PHI_1 Q[7] EN PHI_2 Q[8] VDD VSS DFF_2phase_1
XDFF_2phase_1_3 gc[7] PHI_1 Q[6] EN PHI_2 Q[7] VDD VSS DFF_2phase_1
XDFF_2phase_1_4 gc[6] PHI_1 Q[5] EN PHI_2 Q[6] VDD VSS DFF_2phase_1
XDFF_2phase_1_5 gc[5] PHI_1 Q[4] EN PHI_2 Q[5] VDD VSS DFF_2phase_1
XDFF_2phase_1_6 gc[4] PHI_1 Q[3] EN PHI_2 Q[4] VDD VSS DFF_2phase_1
XDFF_2phase_1_7 gc[3] PHI_1 Q[2] EN PHI_2 Q[3] VDD VSS DFF_2phase_1
XDFF_2phase_1_8 gc[1] PHI_1 D_in EN PHI_2 Q[1] VDD VSS DFF_2phase_1
XDFF_2phase_1_9 gc[2] PHI_1 Q[1] EN PHI_2 Q[2] VDD VSS DFF_2phase_1
.ends

.subckt top vout_s4 vin_s5 vout_s5 vout_lif vin_lif i_in0 vout_0 i_in1 vout_1 i_in2
+ vout_2 i_in3 vout_3 i_in4 vout_4 VAH_bias v_ex v_inh vin_s0 vout_s0 vin_s1 vout_s1
+ vin_s2 vout_s2 vin_s3 vout_s3 vin_s4 enable clk d_in TG_in TG_out TG_clk vss vdd
+ Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
XNO_ClkGen$1_0 TG_clk NO_ClkGen$1_0/phi_2 NO_ClkGen$1_0/phi_1 vdd vss NO_ClkGen$1
XAH_neuron$1_0 vdd i_in3 VAH_bias vout_3 vss AH_neuron$1
XAH_neuron$1_1 vdd i_in2 VAH_bias vout_2 vss AH_neuron$1
XAH_neuron$1_2 vdd i_in1 VAH_bias vout_1 vss AH_neuron$1
XAH_neuron$1_3 vdd i_in0 VAH_bias vout_0 vss AH_neuron$1
Xschmitt_trigger_0 vdd schmitt_trigger_0/out clk vss schmitt_trigger
Xschmitt_trigger_1 vdd schmitt_trigger_1/out d_in vss schmitt_trigger
XTG_bootstrapped_0 NO_ClkGen$1_0/phi_1 vss TG_out NO_ClkGen$1_0/phi_2 TG_in vdd TG_bootstrapped
Xswmatrix_24_by_10_0 vout_lif vin_lif vout_0 i_in0 vout_1 i_in1 vout_2 i_in2 vout_3
+ i_in3 vout_4 i_in4 vout_s5 vin_s5 vout_s4 vin_s4 vout_s3 vout_s1 vin_s3 vout_s2
+ vin_s2 vin_s1 vout_s0 vin_s0 swmatrix_24_by_10_0/D_out schmitt_trigger_0/out schmitt_trigger_1/out
+ swmatrix_24_by_10_0/BUS[1] swmatrix_24_by_10_0/BUS[2] swmatrix_24_by_10_0/BUS[3]
+ swmatrix_24_by_10_0/BUS[4] swmatrix_24_by_10_0/BUS[5] swmatrix_24_by_10_0/BUS[6]
+ swmatrix_24_by_10_0/BUS[7] swmatrix_24_by_10_0/BUS[8] swmatrix_24_by_10_0/BUS[9]
+ swmatrix_24_by_10_0/BUS[10] vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd vdd vdd vdd vdd enable ShiftReg_row_10_2$2_0/PHI_2 ShiftReg_row_10_2$2_0/PHI_1
+ vdd vss vdd vdd swmatrix_24_by_10
Xsynapse_0 v_inh synapse_0/v_ctrl vin_s0 v_ex vdd vout_s0 Q[6] vss synapse
Xsynapse_1 v_inh synapse_1/v_ctrl vin_s1 v_ex vdd vout_s1 Q[5] vss synapse
Xsynapse_2 v_inh synapse_2/v_ctrl vin_s4 v_ex vdd vout_s4 Q[2] vss synapse
Xsynapse_3 v_inh synapse_3/v_ctrl vin_s5 v_ex vdd vout_s5 Q[1] vss synapse
XAH_neuron_0 vdd i_in4 VAH_bias vout_4 vss AH_neuron
XLIF_comp_0 vin_lif Q[7] vout_lif vdd vss LIF_comp
Xsynapse_4 v_inh synapse_4/v_ctrl vin_s2 v_ex vdd vout_s2 Q[4] vss synapse
Xsynapse_5 v_inh synapse_5/v_ctrl vin_s3 v_ex vdd vout_s3 Q[3] vss synapse
XShiftReg_row_10_2$2_0 ShiftReg_row_10_2$2_0/gc[1] ShiftReg_row_10_2$2_0/gc[2] ShiftReg_row_10_2$2_0/gc[3]
+ ShiftReg_row_10_2$2_0/gc[4] ShiftReg_row_10_2$2_0/gc[5] ShiftReg_row_10_2$2_0/gc[6]
+ ShiftReg_row_10_2$2_0/gc[7] ShiftReg_row_10_2$2_0/gc[8] ShiftReg_row_10_2$2_0/gc[9]
+ ShiftReg_row_10_2$2_0/gc[10] ShiftReg_row_10_2$2_0/Q[10] ShiftReg_row_10_2$2_0/PHI_2
+ Q[4] ShiftReg_row_10_2$2_0/Q[9] Q[3] ShiftReg_row_10_2$2_0/Q[8] Q[5] Q[7] Q[6] Q[1]
+ Q[2] enable swmatrix_24_by_10_0/D_out ShiftReg_row_10_2$2_0/PHI_1 vdd vss ShiftReg_row_10_2$2
.ends

