* Extracted by KLayout with GF180MCU LVS runset on : 20/10/2025 01:55

.SUBCKT swmatrix_row_10 E|PHI_1 E|PHI_2 VDD I|ZN|gated_control|gc[1] ZN
+ I|ZN|gated_control|gc[2] I|ZN|gated_control|gc[3] I|ZN|gated_control|gc[4]
+ I|ZN|gated_control|gc[5] I|ZN|gated_control|gc[6] I|ZN|gated_control|gc[7]
+ I|ZN|gated_control|gc[8] I|ZN|gated_control|gc[9] I|ZN|gated_control|gc[10]
+ BUS[1]|T2 BUS[2]|T2 BUS[3]|T2 BUS[4]|T2 BUS[5]|T2 BUS[6]|T2 BUS[7]|T2
+ BUS[8]|T2 BUS[9]|T2 BUS[10]|T2 T1|pin VSS|vss D|Q A1|EN I|ZN A2|D|Q|Q[2]
+ A2|D|Q|Q[3] A2|D|Q|Q[4] A2|D|Q|Q[5] A2|D|Q|Q[6] A2|D|Q|Q[7] A2|D|Q|Q[8]
+ A2|Q|Q[10]|d_out D|D_in A2|D|Q|Q[1] A2|D|Q|Q[9] vss
M$1 T1|pin ZN BUS[1]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$18 T1|pin ZN BUS[2]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$35 T1|pin ZN BUS[3]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$52 T1|pin ZN BUS[4]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$69 T1|pin ZN BUS[5]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$86 T1|pin ZN BUS[6]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$103 T1|pin ZN BUS[7]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$120 T1|pin ZN BUS[8]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$137 T1|pin ZN BUS[9]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$154 T1|pin ZN BUS[10]|T2 VDD pfet_03v3 L=0.28U W=68U AS=19.24P AD=19.24P
+ PS=81.62U PD=81.62U
M$171 VDD I|ZN|gated_control|gc[1] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$172 VDD I|ZN|gated_control|gc[2] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$173 VDD I|ZN|gated_control|gc[3] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$174 VDD I|ZN|gated_control|gc[4] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$175 VDD I|ZN|gated_control|gc[5] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$176 VDD I|ZN|gated_control|gc[6] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$177 VDD I|ZN|gated_control|gc[7] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$178 VDD I|ZN|gated_control|gc[8] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$179 VDD I|ZN|gated_control|gc[9] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$180 VDD I|ZN|gated_control|gc[10] ZN VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$181 VDD E|PHI_1 \$116 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$182 \$117 \$116 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$183 VDD \$183 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$184 VDD E|PHI_2 \$119 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$185 \$120 \$119 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$186 VDD \$185 A2|D|Q|Q[1] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$187 I|ZN A2|D|Q|Q[1] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$188 VDD A1|EN I|ZN VDD pfet_05v0 L=0.5U W=16.45U AS=4.277P AD=7.238P
+ PS=21.65U PD=41.7U
M$189 I|ZN|gated_control|gc[1] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$190 VDD E|PHI_1 \$123 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$191 \$124 \$123 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$192 VDD \$188 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$193 VDD E|PHI_2 \$126 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$194 \$127 \$126 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$195 VDD \$190 A2|D|Q|Q[2] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$196 I|ZN A2|D|Q|Q[2] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$198 I|ZN|gated_control|gc[2] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$199 VDD E|PHI_1 \$130 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$200 \$131 \$130 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$201 VDD \$192 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$202 VDD E|PHI_2 \$133 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$203 \$134 \$133 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$204 VDD \$194 A2|D|Q|Q[3] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$205 I|ZN A2|D|Q|Q[3] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$207 I|ZN|gated_control|gc[3] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$208 VDD E|PHI_1 \$137 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$209 \$138 \$137 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$210 VDD \$196 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$211 VDD E|PHI_2 \$139 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$212 \$140 \$139 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$213 VDD \$199 A2|D|Q|Q[4] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$214 I|ZN A2|D|Q|Q[4] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$216 I|ZN|gated_control|gc[4] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$217 VDD E|PHI_1 \$143 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$218 \$144 \$143 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$219 VDD \$201 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$220 VDD E|PHI_2 \$145 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$221 \$146 \$145 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$222 VDD \$204 A2|D|Q|Q[5] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$223 I|ZN A2|D|Q|Q[5] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$225 I|ZN|gated_control|gc[5] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$226 VDD E|PHI_1 \$149 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$227 \$150 \$149 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$228 VDD \$206 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$229 VDD E|PHI_2 \$152 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$230 \$153 \$152 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$231 VDD \$208 A2|D|Q|Q[6] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$232 I|ZN A2|D|Q|Q[6] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$234 I|ZN|gated_control|gc[6] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$235 VDD E|PHI_1 \$156 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$236 \$157 \$156 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$237 VDD \$210 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$238 VDD E|PHI_2 \$158 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$239 \$159 \$158 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$240 VDD \$213 A2|D|Q|Q[7] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$241 I|ZN A2|D|Q|Q[7] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$243 I|ZN|gated_control|gc[7] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$244 VDD E|PHI_1 \$162 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$245 \$163 \$162 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$246 VDD \$215 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$247 VDD E|PHI_2 \$165 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$248 \$166 \$165 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$249 VDD \$217 A2|D|Q|Q[8] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$250 I|ZN A2|D|Q|Q[8] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$252 I|ZN|gated_control|gc[8] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$253 VDD E|PHI_1 \$169 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$254 \$170 \$169 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$255 VDD \$219 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$256 VDD E|PHI_2 \$172 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$257 \$173 \$172 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$258 VDD \$221 A2|D|Q|Q[9] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$259 I|ZN A2|D|Q|Q[9] VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P AD=0.4277P
+ PS=4.17U PD=2.165U
M$261 I|ZN|gated_control|gc[9] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$262 VDD E|PHI_1 \$175 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$263 \$176 \$175 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$264 VDD \$224 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$265 VDD E|PHI_2 \$178 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$266 \$179 \$178 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$267 VDD \$226 A2|Q|Q[10]|d_out VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P
+ AD=0.8052P PS=4.54U PD=4.54U
M$268 I|ZN A2|Q|Q[10]|d_out VDD VDD pfet_05v0 L=0.5U W=1.645U AS=0.7238P
+ AD=0.4277P PS=4.17U PD=2.165U
M$270 I|ZN|gated_control|gc[10] I|ZN VDD VDD pfet_05v0 L=0.5U W=1.83U
+ AS=0.8052P AD=0.8052P PS=4.54U PD=4.54U
M$271 \$419 D|D_in VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$272 \$183 \$116 \$419 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$273 \$183 \$117 \$421 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$274 VDD \$184 \$421 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$275 \$184 \$183 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$276 \$424 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$277 \$185 \$119 \$424 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$278 \$185 \$120 \$427 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$279 VDD \$186 \$427 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$280 \$186 \$185 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$281 \$433 A2|D|Q|Q[1] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$282 \$188 \$123 \$433 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$283 \$188 \$124 \$436 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$284 VDD \$189 \$436 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$285 \$189 \$188 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$286 \$439 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$287 \$190 \$126 \$439 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$288 \$190 \$127 \$441 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$289 VDD \$191 \$441 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$290 \$191 \$190 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$291 \$447 A2|D|Q|Q[2] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$292 \$192 \$130 \$447 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$293 \$192 \$131 \$449 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$294 VDD \$193 \$449 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$295 \$193 \$192 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$296 \$454 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$297 \$194 \$133 \$454 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$298 \$194 \$134 \$456 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$299 VDD \$195 \$456 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$300 \$195 \$194 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$301 \$461 A2|D|Q|Q[3] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$302 \$196 \$137 \$461 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$303 \$196 \$138 \$464 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$304 VDD \$197 \$464 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$305 \$197 \$196 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$306 \$469 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$307 \$199 \$139 \$469 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$308 \$199 \$140 \$467 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$309 VDD \$200 \$467 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$310 \$200 \$199 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$311 \$475 A2|D|Q|Q[4] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$312 \$201 \$143 \$475 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$313 \$201 \$144 \$477 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$314 VDD \$202 \$477 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$315 \$202 \$201 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$316 \$483 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$317 \$204 \$145 \$483 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$318 \$204 \$146 \$481 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$319 VDD \$205 \$481 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$320 \$205 \$204 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$321 \$489 A2|D|Q|Q[5] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$322 \$206 \$149 \$489 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$323 \$206 \$150 \$492 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$324 VDD \$207 \$492 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$325 \$207 \$206 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$326 \$495 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$327 \$208 \$152 \$495 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$328 \$208 \$153 \$498 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$329 VDD \$209 \$498 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$330 \$209 \$208 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$331 \$503 A2|D|Q|Q[6] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$332 \$210 \$156 \$503 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$333 \$210 \$157 \$506 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$334 VDD \$211 \$506 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$335 \$211 \$210 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$336 \$510 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$337 \$213 \$158 \$510 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$338 \$213 \$159 \$512 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$339 VDD \$214 \$512 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$340 \$214 \$213 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$341 \$517 A2|D|Q|Q[7] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$342 \$215 \$162 \$517 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$343 \$215 \$163 \$520 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$344 VDD \$216 \$520 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$345 \$216 \$215 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$346 \$524 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$347 \$217 \$165 \$524 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$348 \$217 \$166 \$526 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$349 VDD \$218 \$526 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$350 \$218 \$217 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$351 \$531 A2|D|Q|Q[8] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$352 \$219 \$169 \$531 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$353 \$219 \$170 \$534 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$354 VDD \$220 \$534 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$355 \$220 \$219 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$356 \$539 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$357 \$221 \$172 \$539 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$358 \$221 \$173 \$537 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$359 VDD \$222 \$537 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$360 \$222 \$221 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$361 \$546 A2|D|Q|Q[9] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$362 \$224 \$175 \$546 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$363 \$224 \$176 \$548 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$364 VDD \$225 \$548 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$365 \$225 \$224 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$366 \$552 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$367 \$226 \$178 \$552 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$368 \$226 \$179 \$554 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$369 VDD \$227 \$554 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$370 \$227 \$226 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$371 BUS[1]|T2 I|ZN|gated_control|gc[1] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$377 BUS[2]|T2 I|ZN|gated_control|gc[2] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$383 BUS[3]|T2 I|ZN|gated_control|gc[3] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$389 BUS[4]|T2 I|ZN|gated_control|gc[4] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$395 BUS[5]|T2 I|ZN|gated_control|gc[5] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$401 BUS[6]|T2 I|ZN|gated_control|gc[6] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$407 BUS[7]|T2 I|ZN|gated_control|gc[7] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$413 BUS[8]|T2 I|ZN|gated_control|gc[8] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$419 BUS[9]|T2 I|ZN|gated_control|gc[9] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$425 BUS[10]|T2 I|ZN|gated_control|gc[10] T1|pin vss nfet_03v3 L=0.28U W=24U
+ AS=7.64P AD=7.64P PS=31.82U PD=31.82U
M$431 VSS|vss I|ZN|gated_control|gc[1] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$432 VSS|vss \$183 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$433 VSS|vss \$185 A2|D|Q|Q[1] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$434 \$245 A2|D|Q|Q[1] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$435 I|ZN A1|EN \$245 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$436 I|ZN|gated_control|gc[1] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$437 VSS|vss I|ZN|gated_control|gc[2] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$438 VSS|vss \$188 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$439 VSS|vss \$190 A2|D|Q|Q[2] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$440 \$265 A2|D|Q|Q[2] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$441 I|ZN A1|EN \$265 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$442 I|ZN|gated_control|gc[2] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$443 VSS|vss I|ZN|gated_control|gc[3] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$444 VSS|vss \$192 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$445 VSS|vss \$194 A2|D|Q|Q[3] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$446 \$286 A2|D|Q|Q[3] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$447 I|ZN A1|EN \$286 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$448 I|ZN|gated_control|gc[3] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$449 VSS|vss I|ZN|gated_control|gc[4] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$450 VSS|vss \$196 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$451 VSS|vss \$199 A2|D|Q|Q[4] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$452 \$306 A2|D|Q|Q[4] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$453 I|ZN A1|EN \$306 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$454 I|ZN|gated_control|gc[4] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$455 VSS|vss I|ZN|gated_control|gc[5] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$456 VSS|vss \$201 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$457 VSS|vss \$204 A2|D|Q|Q[5] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$458 \$328 A2|D|Q|Q[5] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$459 I|ZN A1|EN \$328 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$460 I|ZN|gated_control|gc[5] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$461 VSS|vss I|ZN|gated_control|gc[6] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$462 VSS|vss \$206 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$463 VSS|vss \$208 A2|D|Q|Q[6] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$464 \$350 A2|D|Q|Q[6] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$465 I|ZN A1|EN \$350 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$466 I|ZN|gated_control|gc[6] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$467 VSS|vss I|ZN|gated_control|gc[7] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$468 VSS|vss \$210 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$469 VSS|vss \$213 A2|D|Q|Q[7] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$470 \$368 A2|D|Q|Q[7] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$471 I|ZN A1|EN \$368 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$472 I|ZN|gated_control|gc[7] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$473 VSS|vss I|ZN|gated_control|gc[8] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$474 VSS|vss \$215 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$475 VSS|vss \$217 A2|D|Q|Q[8] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$476 \$383 A2|D|Q|Q[8] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$477 I|ZN A1|EN \$383 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$478 I|ZN|gated_control|gc[8] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$479 VSS|vss I|ZN|gated_control|gc[9] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$480 VSS|vss \$219 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$481 VSS|vss \$221 A2|D|Q|Q[9] vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$482 \$308 A2|D|Q|Q[9] VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$483 I|ZN A1|EN \$308 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$484 I|ZN|gated_control|gc[9] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$485 VSS|vss I|ZN|gated_control|gc[10] ZN vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$486 VSS|vss \$224 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$487 VSS|vss \$226 A2|Q|Q[10]|d_out vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$488 \$244 A2|Q|Q[10]|d_out VSS|vss vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.2112P PS=3.52U PD=1.64U
M$489 I|ZN A1|EN \$244 vss nfet_05v0 L=0.6U W=1.32U AS=0.2112P AD=0.5808P
+ PS=1.64U PD=3.52U
M$490 I|ZN|gated_control|gc[10] I|ZN VSS|vss vss nfet_05v0 L=0.6U W=1.32U
+ AS=0.5808P AD=0.5808P PS=3.52U PD=3.52U
M$491 VSS|vss E|PHI_1 \$116 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$492 \$117 \$116 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$493 \$231 D|D_in VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$494 \$183 \$117 \$231 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$495 \$230 \$116 \$183 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$496 VSS|vss \$184 \$230 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$497 \$184 \$183 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$498 VSS|vss E|PHI_2 \$119 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$499 \$120 \$119 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$500 \$240 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$501 \$185 \$120 \$240 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$502 \$238 \$119 \$185 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$503 VSS|vss \$186 \$238 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$504 \$186 \$185 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$505 VSS|vss E|PHI_1 \$123 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$506 \$124 \$123 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$507 \$251 A2|D|Q|Q[1] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$508 \$188 \$124 \$251 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$509 \$253 \$123 \$188 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$510 VSS|vss \$189 \$253 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$511 \$189 \$188 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$512 VSS|vss E|PHI_2 \$126 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$513 \$127 \$126 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$514 \$260 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$515 \$190 \$127 \$260 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$516 \$259 \$126 \$190 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$517 VSS|vss \$191 \$259 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$518 \$191 \$190 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$519 VSS|vss E|PHI_1 \$130 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$520 \$131 \$130 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$521 \$274 A2|D|Q|Q[2] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$522 \$192 \$131 \$274 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$523 \$272 \$130 \$192 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$524 VSS|vss \$193 \$272 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$525 \$193 \$192 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$526 VSS|vss E|PHI_2 \$133 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$527 \$134 \$133 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$528 \$281 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$529 \$194 \$134 \$281 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$530 \$284 \$133 \$194 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$531 VSS|vss \$195 \$284 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$532 \$195 \$194 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$533 VSS|vss E|PHI_1 \$137 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$534 \$138 \$137 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$535 \$295 A2|D|Q|Q[3] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$536 \$196 \$138 \$295 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$537 \$293 \$137 \$196 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$538 VSS|vss \$197 \$293 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$539 \$197 \$196 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$540 VSS|vss E|PHI_2 \$139 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$541 \$140 \$139 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$542 \$301 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$543 \$199 \$140 \$301 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$544 \$303 \$139 \$199 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$545 VSS|vss \$200 \$303 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$546 \$200 \$199 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$547 VSS|vss E|PHI_1 \$143 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$548 \$144 \$143 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$549 \$314 A2|D|Q|Q[4] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$550 \$201 \$144 \$314 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$551 \$315 \$143 \$201 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$552 VSS|vss \$202 \$315 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$553 \$202 \$201 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$554 VSS|vss E|PHI_2 \$145 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$555 \$146 \$145 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$556 \$322 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$557 \$204 \$146 \$322 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$558 \$321 \$145 \$204 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$559 VSS|vss \$205 \$321 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$560 \$205 \$204 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$561 VSS|vss E|PHI_1 \$149 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$562 \$150 \$149 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$563 \$335 A2|D|Q|Q[5] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$564 \$206 \$150 \$335 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$565 \$336 \$149 \$206 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$566 VSS|vss \$207 \$336 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$567 \$207 \$206 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$568 VSS|vss E|PHI_2 \$152 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$569 \$153 \$152 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$570 \$343 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$571 \$208 \$153 \$343 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$572 \$344 \$152 \$208 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$573 VSS|vss \$209 \$344 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$574 \$209 \$208 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$575 VSS|vss E|PHI_1 \$156 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$576 \$157 \$156 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$577 \$356 A2|D|Q|Q[6] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$578 \$210 \$157 \$356 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$579 \$357 \$156 \$210 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$580 VSS|vss \$211 \$357 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$581 \$211 \$210 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$582 VSS|vss E|PHI_2 \$158 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$583 \$159 \$158 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$584 \$365 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$585 \$213 \$159 \$365 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$586 \$364 \$158 \$213 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$587 VSS|vss \$214 \$364 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$588 \$214 \$213 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$589 VSS|vss E|PHI_1 \$162 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$590 \$163 \$162 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$591 \$377 A2|D|Q|Q[7] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$592 \$215 \$163 \$377 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$593 \$375 \$162 \$215 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$594 VSS|vss \$216 \$375 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$595 \$216 \$215 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$596 VSS|vss E|PHI_2 \$165 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$597 \$166 \$165 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$598 \$385 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$599 \$217 \$166 \$385 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$600 \$384 \$165 \$217 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$601 VSS|vss \$218 \$384 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$602 \$218 \$217 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$603 VSS|vss E|PHI_1 \$169 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$604 \$170 \$169 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$605 \$351 A2|D|Q|Q[8] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$606 \$219 \$170 \$351 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$607 \$347 \$169 \$219 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$608 VSS|vss \$220 \$347 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$609 \$220 \$219 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$610 VSS|vss E|PHI_2 \$172 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$611 \$173 \$172 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$612 \$325 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$613 \$221 \$173 \$325 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$614 \$329 \$172 \$221 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$615 VSS|vss \$222 \$329 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$616 \$222 \$221 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$617 VSS|vss E|PHI_1 \$175 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$618 \$176 \$175 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$619 \$280 A2|D|Q|Q[9] VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$620 \$224 \$176 \$280 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$621 \$283 \$175 \$224 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$622 VSS|vss \$225 \$283 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$623 \$225 \$224 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$624 VSS|vss E|PHI_2 \$178 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$625 \$179 \$178 VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$626 \$257 D|Q VSS|vss vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$627 \$226 \$179 \$257 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$628 \$261 \$178 \$226 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$629 VSS|vss \$227 \$261 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$630 \$227 \$226 VSS|vss vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
.ENDS swmatrix_row_10
