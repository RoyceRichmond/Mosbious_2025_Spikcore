* NGSPICE file created from TG_bootstrapped.ext - technology: gf180mcuD

.subckt TG_bootstrapped_pex vdd vss clk nclk vin vout
X0 vout.t26 a_5673_n171.t4 vin.t27 vss.t17 nfet_03v3 ad=2.38815p pd=9.05u as=1.0179p ps=4.435u w=3.915u l=0.42u
X1 vin.t23 a_5673_n171.t5 vout.t25 vss.t16 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X2 vin.t2 a_5297_1329.t4 vout.t2 vdd.t31 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X3 a_8039_2775# a_5944_2919# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X4 vin.t31 clk.t0 a_8039_2775# vss.t23 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X5 vin.t8 a_5297_1329.t5 vout.t7 vdd.t30 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X6 vout.t4 a_5297_1329.t6 vin.t4 vdd.t29 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X7 vout.t6 a_5297_1329.t7 vin.t7 vdd.t28 pfet_03v3 ad=2.028p pd=7.54u as=0.8112p ps=3.64u w=3.12u l=0.42u
X8 vin.t10 a_5297_1329.t8 vout.t9 vdd.t27 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X9 vin.t1 a_5297_1329.t9 vout.t1 vdd.t26 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X10 vss.t1 nclk.t0 a_5673_n171.t1 vss.t0 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X11 vout.t10 a_5297_1329.t10 vin.t12 vdd.t25 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X12 vin.t3 a_5297_1329.t11 vout.t3 vdd.t24 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X13 vin.t6 a_5297_1329.t12 vout.t5 vdd.t23 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X14 a_8034_n1134# nclk.t1 vss.t20 vss.t19 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X15 vin.t11 nclk.t2 a_8034_n1134# vdd.t5 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X16 vin.t28 a_5673_n171.t6 vout.t24 vss.t15 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X17 vout.t23 a_5673_n171.t7 vin.t26 vss.t14 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X18 a_5944_2919# clk.t1 vss.t26 vss.t25 nfet_03v3 ad=0.3416p pd=2.34u as=0.3416p ps=2.34u w=0.56u l=0.28u
X19 vout.t22 a_5673_n171.t8 vin.t21 vss.t13 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X20 vout.t21 a_5673_n171.t9 vin.t17 vss.t12 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X21 vdd.t11 clk.t2 a_5297_1329.t2 vdd.t10 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X22 vin.t19 a_5673_n171.t10 vout.t20 vss.t11 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X23 a_5939_n1022# clk.t3 vdd.t8 vdd.t7 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X24 a_5297_1329.t0 nclk.t3 a_5944_2919# vdd.t1 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X25 a_5673_n171.t0 nclk.t4 a_5939_n1022# vdd.t0 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X26 vin.t9 a_5297_1329.t13 vout.t8 vdd.t22 pfet_03v3 ad=0.8112p pd=3.64u as=2.028p ps=7.54u w=3.12u l=0.42u
X27 vout.t0 a_5297_1329.t14 vin.t0 vdd.t21 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X28 vout.t27 a_5297_1329.t15 vin.t29 vdd.t20 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X29 vout.t35 a_5297_1329.t16 vin.t39 vdd.t19 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X30 vin.t38 a_5297_1329.t17 vout.t34 vdd.t18 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X31 a_8034_n1134# a_5939_n1022# cap_mim_2f0_m4m5_noshield c_width=7u c_length=8u
X32 vin.t5 nclk.t5 a_8039_2775# vdd.t2 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X33 vdd.t6 nclk.t6 a_5297_1329.t1 vss.t18 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X34 a_5297_1329.t3 clk.t4 a_5944_2919# vss.t27 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X35 vin.t25 a_5673_n171.t11 vout.t19 vss.t10 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X36 vss.t24 clk.t5 a_5673_n171.t3 vdd.t9 pfet_03v3 ad=1.092p pd=4.66u as=1.092p ps=4.66u w=1.68u l=0.84u
X37 vin.t18 a_5673_n171.t12 vout.t18 vss.t9 nfet_03v3 ad=1.0179p pd=4.435u as=2.38815p ps=9.05u w=3.915u l=0.42u
X38 vin.t15 a_5673_n171.t13 vout.t17 vss.t8 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X39 vout.t16 a_5673_n171.t14 vin.t20 vss.t7 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X40 vdd.t4 nclk.t7 a_8039_2775# vdd.t3 pfet_03v3 ad=0.728p pd=3.54u as=0.728p ps=3.54u w=1.12u l=0.28u
X41 vout.t15 a_5673_n171.t15 vin.t13 vss.t6 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X42 vout.t33 a_5297_1329.t18 vin.t37 vdd.t17 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X43 vin.t33 a_5297_1329.t19 vout.t29 vdd.t16 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X44 vout.t32 a_5297_1329.t20 vin.t36 vdd.t15 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X45 vout.t30 a_5297_1329.t21 vin.t34 vdd.t14 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X46 vout.t31 a_5297_1329.t22 vin.t35 vdd.t13 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X47 vin.t32 a_5297_1329.t23 vout.t28 vdd.t12 pfet_03v3 ad=0.8112p pd=3.64u as=0.8112p ps=3.64u w=3.12u l=0.42u
X48 vout.t14 a_5673_n171.t16 vin.t24 vss.t5 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X49 vin.t30 clk.t6 a_8034_n1134# vss.t22 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
X50 vout.t13 a_5673_n171.t17 vin.t22 vss.t4 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X51 vin.t14 a_5673_n171.t18 vout.t12 vss.t3 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X52 vin.t16 a_5673_n171.t19 vout.t11 vss.t2 nfet_03v3 ad=1.0179p pd=4.435u as=1.0179p ps=4.435u w=3.915u l=0.42u
X53 a_5673_n171.t2 clk.t7 a_5939_n1022# vss.t21 nfet_03v3 ad=0.5124p pd=2.9u as=0.5124p ps=2.9u w=0.84u l=0.84u
R0 a_5673_n171.n5 a_5673_n171.t12 50.5346
R1 a_5673_n171.n14 a_5673_n171.t4 50.5346
R2 a_5673_n171.n5 a_5673_n171.t17 50.3231
R3 a_5673_n171.n6 a_5673_n171.t5 50.3231
R4 a_5673_n171.n7 a_5673_n171.t8 50.3231
R5 a_5673_n171.n8 a_5673_n171.t13 50.3231
R6 a_5673_n171.n9 a_5673_n171.t16 50.3231
R7 a_5673_n171.n12 a_5673_n171.t6 50.3231
R8 a_5673_n171.n11 a_5673_n171.t9 50.3231
R9 a_5673_n171.n20 a_5673_n171.t10 50.3231
R10 a_5673_n171.n19 a_5673_n171.t15 50.3231
R11 a_5673_n171.n18 a_5673_n171.t18 50.3231
R12 a_5673_n171.n17 a_5673_n171.t7 50.3231
R13 a_5673_n171.n16 a_5673_n171.t11 50.3231
R14 a_5673_n171.n15 a_5673_n171.t14 50.3231
R15 a_5673_n171.n14 a_5673_n171.t19 50.3231
R16 a_5673_n171.n28 a_5673_n171.t2 9.65132
R17 a_5673_n171.n3 a_5673_n171.t1 9.65118
R18 a_5673_n171.n22 a_5673_n171.n10 9.0005
R19 a_5673_n171.n22 a_5673_n171.n13 9.0005
R20 a_5673_n171.n22 a_5673_n171.n4 9.0005
R21 a_5673_n171.n22 a_5673_n171.n21 9.0005
R22 a_5673_n171.n25 a_5673_n171.n23 4.5005
R23 a_5673_n171.n26 a_5673_n171.n2 4.5005
R24 a_5673_n171.n27 a_5673_n171.n26 4.5005
R25 a_5673_n171.n26 a_5673_n171.n25 4.5005
R26 a_5673_n171.n3 a_5673_n171.t3 3.70851
R27 a_5673_n171.t0 a_5673_n171.n28 3.70835
R28 a_5673_n171.n24 a_5673_n171.n1 2.24455
R29 a_5673_n171.n23 a_5673_n171.n0 2.24204
R30 a_5673_n171.n25 a_5673_n171.n3 1.04078
R31 a_5673_n171.n28 a_5673_n171.n27 1.03838
R32 a_5673_n171.n15 a_5673_n171.n14 0.212
R33 a_5673_n171.n16 a_5673_n171.n15 0.212
R34 a_5673_n171.n17 a_5673_n171.n16 0.212
R35 a_5673_n171.n18 a_5673_n171.n17 0.212
R36 a_5673_n171.n19 a_5673_n171.n18 0.212
R37 a_5673_n171.n9 a_5673_n171.n8 0.212
R38 a_5673_n171.n8 a_5673_n171.n7 0.212
R39 a_5673_n171.n7 a_5673_n171.n6 0.212
R40 a_5673_n171.n6 a_5673_n171.n5 0.212
R41 a_5673_n171.n21 a_5673_n171.n20 0.147875
R42 a_5673_n171.n11 a_5673_n171.n4 0.134375
R43 a_5673_n171.n23 a_5673_n171.n22 0.122181
R44 a_5673_n171.n13 a_5673_n171.n12 0.120875
R45 a_5673_n171.n10 a_5673_n171.n9 0.107375
R46 a_5673_n171.n12 a_5673_n171.n10 0.105125
R47 a_5673_n171.n13 a_5673_n171.n11 0.091625
R48 a_5673_n171.n20 a_5673_n171.n4 0.078125
R49 a_5673_n171.n21 a_5673_n171.n19 0.064625
R50 a_5673_n171.n25 a_5673_n171.n24 0.0365
R51 a_5673_n171.n24 a_5673_n171.n2 0.0365
R52 a_5673_n171.n27 a_5673_n171.n0 0.0189283
R53 a_5673_n171.n2 a_5673_n171.n0 0.0189283
R54 a_5673_n171.n26 a_5673_n171.n1 0.013894
R55 a_5673_n171.n23 a_5673_n171.n1 0.013894
R56 vin.n24 vin.t31 18.882
R57 vin.n26 vin.n25 10.1447
R58 vin.n25 vin.t30 9.92542
R59 vin.n24 vin.t5 7.98552
R60 vin.n25 vin.t11 3.48383
R61 vin.n22 vin.n20 2.12064
R62 vin.n80 vin.n78 2.12064
R63 vin.n22 vin.n21 2.05296
R64 vin.n36 vin.n35 2.05296
R65 vin.n16 vin.n15 2.05296
R66 vin.n51 vin.n50 2.05296
R67 vin.n10 vin.n9 2.05296
R68 vin.n65 vin.n64 2.05296
R69 vin.n4 vin.n3 2.05296
R70 vin.n80 vin.n79 2.05296
R71 vin.n29 vin.n28 1.87421
R72 vin.n2 vin.n1 1.86774
R73 vin.n31 vin.n30 1.86521
R74 vin.n44 vin.n43 1.86521
R75 vin.n13 vin.n12 1.86521
R76 vin.n58 vin.n57 1.86521
R77 vin.n7 vin.n6 1.86521
R78 vin.n72 vin.n71 1.86521
R79 vin.n82 vin.n81 1.5005
R80 vin.n77 vin.n0 1.5005
R81 vin.n76 vin.n75 1.5005
R82 vin.n66 vin.n5 1.5005
R83 vin.n68 vin.n67 1.5005
R84 vin.n63 vin.n8 1.5005
R85 vin.n62 vin.n61 1.5005
R86 vin.n52 vin.n11 1.5005
R87 vin.n54 vin.n53 1.5005
R88 vin.n49 vin.n14 1.5005
R89 vin.n48 vin.n47 1.5005
R90 vin.n38 vin.n17 1.5005
R91 vin.n40 vin.n39 1.5005
R92 vin.n37 vin.n19 1.5005
R93 vin.n34 vin.n33 1.5005
R94 vin.n27 vin.n23 1.5005
R95 vin.n26 vin.n24 1.13439
R96 vin.n82 vin.n2 1.1255
R97 vin.n73 vin.n0 1.1255
R98 vin.n75 vin.n74 1.1255
R99 vin.n70 vin.n5 1.1255
R100 vin.n69 vin.n68 1.1255
R101 vin.n59 vin.n8 1.1255
R102 vin.n61 vin.n60 1.1255
R103 vin.n56 vin.n11 1.1255
R104 vin.n55 vin.n54 1.1255
R105 vin.n45 vin.n14 1.1255
R106 vin.n47 vin.n46 1.1255
R107 vin.n42 vin.n17 1.1255
R108 vin.n41 vin.n40 1.1255
R109 vin.n19 vin.n18 1.1255
R110 vin.n33 vin.n32 1.1255
R111 vin.n29 vin.n27 1.1255
R112 vin vin.n82 0.601237
R113 vin.n78 vin.t36 0.583833
R114 vin.n78 vin.t9 0.583833
R115 vin.n79 vin.t0 0.583833
R116 vin.n79 vin.t8 0.583833
R117 vin.n3 vin.t12 0.583833
R118 vin.n3 vin.t32 0.583833
R119 vin.n64 vin.t34 0.583833
R120 vin.n64 vin.t38 0.583833
R121 vin.n9 vin.t29 0.583833
R122 vin.n9 vin.t10 0.583833
R123 vin.n50 vin.t39 0.583833
R124 vin.n50 vin.t1 0.583833
R125 vin.n15 vin.t4 0.583833
R126 vin.n15 vin.t33 0.583833
R127 vin.n35 vin.t35 0.583833
R128 vin.n35 vin.t3 0.583833
R129 vin.n21 vin.t37 0.583833
R130 vin.n21 vin.t6 0.583833
R131 vin.n20 vin.t7 0.583833
R132 vin.n20 vin.t2 0.583833
R133 vin.n1 vin.t22 0.418891
R134 vin.n1 vin.t18 0.418891
R135 vin.n71 vin.t21 0.418891
R136 vin.n71 vin.t23 0.418891
R137 vin.n6 vin.t24 0.418891
R138 vin.n6 vin.t15 0.418891
R139 vin.n57 vin.t17 0.418891
R140 vin.n57 vin.t28 0.418891
R141 vin.n12 vin.t13 0.418891
R142 vin.n12 vin.t19 0.418891
R143 vin.n43 vin.t26 0.418891
R144 vin.n43 vin.t14 0.418891
R145 vin.n30 vin.t20 0.418891
R146 vin.n30 vin.t25 0.418891
R147 vin.n28 vin.t27 0.418891
R148 vin.n28 vin.t16 0.418891
R149 vin.n34 vin.n23 0.0311
R150 vin.n39 vin.n37 0.0311
R151 vin.n39 vin.n38 0.0311
R152 vin.n49 vin.n48 0.0311
R153 vin.n53 vin.n52 0.0311
R154 vin.n63 vin.n62 0.0311
R155 vin.n67 vin.n66 0.0311
R156 vin.n77 vin.n76 0.0311
R157 vin.n81 vin.n77 0.0311
R158 vin.n48 vin.n16 0.02966
R159 vin.n66 vin.n4 0.02786
R160 vin.n36 vin.n34 0.02606
R161 vin.n32 vin.n29 0.0244062
R162 vin.n41 vin.n18 0.0244062
R163 vin.n42 vin.n41 0.0244062
R164 vin.n46 vin.n45 0.0244062
R165 vin.n56 vin.n55 0.0244062
R166 vin.n60 vin.n59 0.0244062
R167 vin.n70 vin.n69 0.0244062
R168 vin.n74 vin.n73 0.0244062
R169 vin.n73 vin.n2 0.0244062
R170 vin.n46 vin.n44 0.0232812
R171 vin.n53 vin.n51 0.02318
R172 vin.n72 vin.n70 0.021875
R173 vin.n65 vin.n63 0.02138
R174 vin.n32 vin.n31 0.0204687
R175 vin.n55 vin.n13 0.0182187
R176 vin.n59 vin.n7 0.0168125
R177 vin.n62 vin.n10 0.0167
R178 vin.n52 vin.n10 0.0149
R179 vin.n60 vin.n58 0.0131563
R180 vin.n23 vin.n22 0.01202
R181 vin.n58 vin.n56 0.01175
R182 vin.n67 vin.n65 0.01022
R183 vin.n33 vin.n27 0.0084729
R184 vin.n33 vin.n19 0.0084729
R185 vin.n40 vin.n19 0.0084729
R186 vin.n40 vin.n17 0.0084729
R187 vin.n47 vin.n17 0.0084729
R188 vin.n47 vin.n14 0.0084729
R189 vin.n54 vin.n14 0.0084729
R190 vin.n54 vin.n11 0.0084729
R191 vin.n61 vin.n11 0.0084729
R192 vin.n61 vin.n8 0.0084729
R193 vin.n68 vin.n8 0.0084729
R194 vin.n68 vin.n5 0.0084729
R195 vin.n75 vin.n5 0.0084729
R196 vin.n75 vin.n0 0.0084729
R197 vin.n82 vin.n0 0.0084729
R198 vin.n51 vin.n49 0.00842
R199 vin.n69 vin.n7 0.00809375
R200 vin.n45 vin.n13 0.0066875
R201 vin.n37 vin.n36 0.00554
R202 vin.n31 vin.n18 0.0044375
R203 vin.n76 vin.n4 0.00374
R204 vin.n81 vin.n80 0.00374
R205 vin.n74 vin.n72 0.00303125
R206 vin.n27 vin.n26 0.00218838
R207 vin.n38 vin.n16 0.00194
R208 vin.n44 vin.n42 0.001625
R209 vout.n1 vout.t6 2.56303
R210 vout.n28 vout.t8 2.56303
R211 vout.n29 vout.n26 2.31025
R212 vout.n31 vout.n26 2.2505
R213 vout.n33 vout.n32 2.2505
R214 vout.n35 vout.n34 2.2505
R215 vout.n36 vout.n20 2.2505
R216 vout.n39 vout.n38 2.2505
R217 vout.n40 vout.n19 2.2505
R218 vout.n42 vout.n41 2.2505
R219 vout.n44 vout.n16 2.2505
R220 vout.n46 vout.n45 2.2505
R221 vout.n48 vout.n47 2.2505
R222 vout.n49 vout.n10 2.2505
R223 vout.n52 vout.n51 2.2505
R224 vout.n53 vout.n9 2.2505
R225 vout.n55 vout.n54 2.2505
R226 vout.n57 vout.n6 2.2505
R227 vout.n59 vout.n58 2.2505
R228 vout.n61 vout.n60 2.2505
R229 vout.n62 vout.n0 2.2505
R230 vout.n65 vout.n64 2.2505
R231 vout.n28 vout.t18 2.24523
R232 vout.n1 vout.t26 2.24523
R233 vout.n5 vout.n4 1.60155
R234 vout.n56 vout.n8 1.60155
R235 vout.n50 vout.n12 1.60155
R236 vout.n15 vout.n14 1.60155
R237 vout.n43 vout.n18 1.60155
R238 vout.n37 vout.n22 1.60155
R239 vout.n25 vout.n24 1.60155
R240 vout.n63 vout.n2 1.47822
R241 vout.n5 vout.n3 1.47822
R242 vout.n56 vout.n7 1.47822
R243 vout.n50 vout.n11 1.47822
R244 vout.n15 vout.n13 1.47822
R245 vout.n43 vout.n17 1.47822
R246 vout.n37 vout.n21 1.47822
R247 vout.n25 vout.n23 1.47822
R248 vout.n30 vout.n27 1.47822
R249 vout vout.n65 1.02411
R250 vout.n2 vout.t2 0.583833
R251 vout.n2 vout.t33 0.583833
R252 vout.n3 vout.t5 0.583833
R253 vout.n3 vout.t31 0.583833
R254 vout.n7 vout.t3 0.583833
R255 vout.n7 vout.t4 0.583833
R256 vout.n11 vout.t29 0.583833
R257 vout.n11 vout.t35 0.583833
R258 vout.n13 vout.t1 0.583833
R259 vout.n13 vout.t27 0.583833
R260 vout.n17 vout.t9 0.583833
R261 vout.n17 vout.t30 0.583833
R262 vout.n21 vout.t34 0.583833
R263 vout.n21 vout.t10 0.583833
R264 vout.n23 vout.t28 0.583833
R265 vout.n23 vout.t0 0.583833
R266 vout.n27 vout.t7 0.583833
R267 vout.n27 vout.t32 0.583833
R268 vout.n4 vout.t11 0.418891
R269 vout.n4 vout.t16 0.418891
R270 vout.n8 vout.t19 0.418891
R271 vout.n8 vout.t23 0.418891
R272 vout.n12 vout.t12 0.418891
R273 vout.n12 vout.t15 0.418891
R274 vout.n14 vout.t20 0.418891
R275 vout.n14 vout.t21 0.418891
R276 vout.n18 vout.t24 0.418891
R277 vout.n18 vout.t14 0.418891
R278 vout.n22 vout.t17 0.418891
R279 vout.n22 vout.t22 0.418891
R280 vout.n24 vout.t25 0.418891
R281 vout.n24 vout.t13 0.418891
R282 vout.n62 vout.n61 0.0605
R283 vout.n58 vout.n57 0.0605
R284 vout.n55 vout.n9 0.0605
R285 vout.n51 vout.n9 0.0605
R286 vout.n49 vout.n48 0.0605
R287 vout.n45 vout.n44 0.0605
R288 vout.n42 vout.n19 0.0605
R289 vout.n38 vout.n19 0.0605
R290 vout.n36 vout.n35 0.0605
R291 vout.n32 vout.n31 0.0605
R292 vout.n65 vout.n0 0.060251
R293 vout.n60 vout.n0 0.060251
R294 vout.n60 vout.n59 0.060251
R295 vout.n59 vout.n6 0.060251
R296 vout.n54 vout.n6 0.060251
R297 vout.n54 vout.n53 0.060251
R298 vout.n53 vout.n52 0.060251
R299 vout.n52 vout.n10 0.060251
R300 vout.n47 vout.n10 0.060251
R301 vout.n47 vout.n46 0.060251
R302 vout.n46 vout.n16 0.060251
R303 vout.n41 vout.n16 0.060251
R304 vout.n41 vout.n40 0.060251
R305 vout.n40 vout.n39 0.060251
R306 vout.n39 vout.n20 0.060251
R307 vout.n34 vout.n20 0.060251
R308 vout.n34 vout.n33 0.060251
R309 vout.n33 vout.n26 0.060251
R310 vout.n63 vout.n62 0.05525
R311 vout.n31 vout.n30 0.05375
R312 vout.n50 vout.n49 0.05225
R313 vout.n44 vout.n43 0.05075
R314 vout.n37 vout.n36 0.04925
R315 vout.n57 vout.n56 0.04775
R316 vout.n58 vout.n5 0.03425
R317 vout.n35 vout.n25 0.03275
R318 vout.n45 vout.n15 0.03125
R319 vout.n48 vout.n15 0.02975
R320 vout.n32 vout.n25 0.02825
R321 vout.n61 vout.n5 0.02675
R322 vout.n56 vout.n55 0.01325
R323 vout.n38 vout.n37 0.01175
R324 vout.n43 vout.n42 0.01025
R325 vout.n51 vout.n50 0.00875
R326 vout.n30 vout.n29 0.00725
R327 vout.n64 vout.n1 0.00575
R328 vout.n64 vout.n63 0.00575
R329 vout.n29 vout.n28 0.00425
R330 vss.n15 vss.n5 21125
R331 vss.n24 vss.t21 5432.3
R332 vss.n25 vss.n24 4678.74
R333 vss.n15 vss.n14 3658.85
R334 vss.t19 vss.n15 2578.99
R335 vss.t22 vss.t0 1060.25
R336 vss.t18 vss.t23 920.038
R337 vss.n23 vss.t0 480.928
R338 vss.t21 vss.n23 480.928
R339 vss.n20 vss.t22 470.882
R340 vss.t27 vss.n5 467.32
R341 vss.n24 vss.t9 418.368
R342 vss.n7 vss.t18 416.243
R343 vss.n7 vss.t27 416.243
R344 vss.n14 vss.t23 406.25
R345 vss.n19 vss.t17 358.844
R346 vss.t17 vss.t2 319.728
R347 vss.t2 vss.t7 319.728
R348 vss.t7 vss.t10 319.728
R349 vss.t10 vss.t14 319.728
R350 vss.t14 vss.t3 319.728
R351 vss.t3 vss.t6 319.728
R352 vss.t6 vss.t11 319.728
R353 vss.t11 vss.t12 319.728
R354 vss.t12 vss.t15 319.728
R355 vss.t15 vss.t5 319.728
R356 vss.t5 vss.t8 319.728
R357 vss.t8 vss.t13 319.728
R358 vss.t13 vss.t16 319.728
R359 vss.t16 vss.t4 319.728
R360 vss.t4 vss.t9 319.728
R361 vss.n20 vss.n19 301.611
R362 vss.n5 vss.t25 267.625
R363 vss.n25 vss.t25 229.131
R364 vss.n16 vss.t19 175.298
R365 vss.n18 vss.n16 86.9476
R366 vss.n19 vss.n18 37.1634
R367 vss.n14 vss.n13 19.8888
R368 vss.n21 vss.n20 19.6851
R369 vss.n4 vss.t20 10.877
R370 vss.n26 vss.t26 10.8546
R371 vss.n16 vss.n4 10.4837
R372 vss.n26 vss.n25 10.4462
R373 vss.n2 vss.t1 9.6559
R374 vss.n21 vss.n4 9.22213
R375 vss.n27 vss.n26 7.16341
R376 vss.n9 vss.n0 4.59325
R377 vss.n11 vss.n8 4.5005
R378 vss.n10 vss.n6 4.5005
R379 vss.n12 vss.n11 4.5005
R380 vss.n18 vss.n17 3.80854
R381 vss.n2 vss.t24 3.71674
R382 vss.n23 vss.n22 3.37699
R383 vss.n3 vss.n2 2.94978
R384 vss.n9 vss.n8 2.20487
R385 vss.n17 vss.n3 1.34213
R386 vss.n22 vss.n1 1.02307
R387 vss.n13 vss.n1 0.918196
R388 vss.n22 vss.n21 0.4415
R389 vss vss.n27 0.359439
R390 vss.n8 vss.n7 0.298561
R391 vss.n13 vss.n12 0.280052
R392 vss.n27 vss.n0 0.244392
R393 vss.n17 vss.n1 0.201851
R394 vss.n11 vss.n10 0.188872
R395 vss.n21 vss.n3 0.176
R396 vss.n10 vss.n9 0.0932551
R397 vss.n12 vss.n6 0.0387075
R398 vss.n6 vss.n0 0.0387075
R399 a_5297_1329.n3 a_5297_1329.t13 43.8541
R400 a_5297_1329.n14 a_5297_1329.t7 43.8541
R401 a_5297_1329.n3 a_5297_1329.t20 43.6315
R402 a_5297_1329.n4 a_5297_1329.t5 43.6315
R403 a_5297_1329.n5 a_5297_1329.t14 43.6315
R404 a_5297_1329.n6 a_5297_1329.t23 43.6315
R405 a_5297_1329.n7 a_5297_1329.t10 43.6315
R406 a_5297_1329.n8 a_5297_1329.t17 43.6315
R407 a_5297_1329.n9 a_5297_1329.t21 43.6315
R408 a_5297_1329.n12 a_5297_1329.t8 43.6315
R409 a_5297_1329.n11 a_5297_1329.t15 43.6315
R410 a_5297_1329.n22 a_5297_1329.t9 43.6315
R411 a_5297_1329.n21 a_5297_1329.t16 43.6315
R412 a_5297_1329.n20 a_5297_1329.t19 43.6315
R413 a_5297_1329.n19 a_5297_1329.t6 43.6315
R414 a_5297_1329.n18 a_5297_1329.t11 43.6315
R415 a_5297_1329.n17 a_5297_1329.t22 43.6315
R416 a_5297_1329.n16 a_5297_1329.t12 43.6315
R417 a_5297_1329.n15 a_5297_1329.t18 43.6315
R418 a_5297_1329.n14 a_5297_1329.t4 43.6315
R419 a_5297_1329.n26 a_5297_1329.t1 9.65161
R420 a_5297_1329.n32 a_5297_1329.t3 9.65118
R421 a_5297_1329.n24 a_5297_1329.n10 9.0005
R422 a_5297_1329.n24 a_5297_1329.n13 9.0005
R423 a_5297_1329.n24 a_5297_1329.n2 9.0005
R424 a_5297_1329.n24 a_5297_1329.n23 9.0005
R425 a_5297_1329.n29 a_5297_1329.n27 4.5005
R426 a_5297_1329.n30 a_5297_1329.n25 4.5005
R427 a_5297_1329.n31 a_5297_1329.n30 4.5005
R428 a_5297_1329.n30 a_5297_1329.n29 4.5005
R429 a_5297_1329.t0 a_5297_1329.n32 3.70851
R430 a_5297_1329.n26 a_5297_1329.t2 3.7081
R431 a_5297_1329.n28 a_5297_1329.n1 2.24497
R432 a_5297_1329.n27 a_5297_1329.n0 2.24204
R433 a_5297_1329.n29 a_5297_1329.n26 1.04096
R434 a_5297_1329.n32 a_5297_1329.n31 1.03826
R435 a_5297_1329.n9 a_5297_1329.n8 0.223132
R436 a_5297_1329.n8 a_5297_1329.n7 0.223132
R437 a_5297_1329.n7 a_5297_1329.n6 0.223132
R438 a_5297_1329.n6 a_5297_1329.n5 0.223132
R439 a_5297_1329.n5 a_5297_1329.n4 0.223132
R440 a_5297_1329.n4 a_5297_1329.n3 0.223132
R441 a_5297_1329.n15 a_5297_1329.n14 0.223132
R442 a_5297_1329.n16 a_5297_1329.n15 0.223132
R443 a_5297_1329.n17 a_5297_1329.n16 0.223132
R444 a_5297_1329.n18 a_5297_1329.n17 0.223132
R445 a_5297_1329.n19 a_5297_1329.n18 0.223132
R446 a_5297_1329.n20 a_5297_1329.n19 0.223132
R447 a_5297_1329.n21 a_5297_1329.n20 0.223132
R448 a_5297_1329.n23 a_5297_1329.n22 0.153263
R449 a_5297_1329.n11 a_5297_1329.n2 0.139053
R450 a_5297_1329.n13 a_5297_1329.n12 0.124842
R451 a_5297_1329.n30 a_5297_1329.n24 0.114452
R452 a_5297_1329.n10 a_5297_1329.n9 0.110632
R453 a_5297_1329.n12 a_5297_1329.n10 0.108263
R454 a_5297_1329.n13 a_5297_1329.n11 0.0940526
R455 a_5297_1329.n22 a_5297_1329.n2 0.0798421
R456 a_5297_1329.n23 a_5297_1329.n21 0.0656316
R457 a_5297_1329.n29 a_5297_1329.n28 0.0365
R458 a_5297_1329.n28 a_5297_1329.n25 0.0365
R459 a_5297_1329.n31 a_5297_1329.n0 0.0189283
R460 a_5297_1329.n25 a_5297_1329.n0 0.0189283
R461 a_5297_1329.n30 a_5297_1329.n1 0.0130643
R462 a_5297_1329.n27 a_5297_1329.n1 0.0130643
R463 vdd.t0 vdd.t7 1167.16
R464 vdd.t10 vdd.t2 1138.89
R465 vdd.t5 vdd.t9 1132.35
R466 vdd.n1 vdd.t3 888.654
R467 vdd.n10 vdd.t5 522.399
R468 vdd.t3 vdd.n0 522.338
R469 vdd.t7 vdd.n8 522.322
R470 vdd.n3 vdd.t10 517.273
R471 vdd.n3 vdd.t1 517.273
R472 vdd.t9 vdd.n9 517.273
R473 vdd.n9 vdd.t0 517.273
R474 vdd.t2 vdd.n1 513.072
R475 vdd.n11 vdd.t28 304.387
R476 vdd.t28 vdd.t31 208.889
R477 vdd.t31 vdd.t17 208.889
R478 vdd.t17 vdd.t23 208.889
R479 vdd.t23 vdd.t13 208.889
R480 vdd.t13 vdd.t24 208.889
R481 vdd.t24 vdd.t29 208.889
R482 vdd.t29 vdd.t16 208.889
R483 vdd.t16 vdd.t19 208.889
R484 vdd.t19 vdd.t26 208.889
R485 vdd.t26 vdd.t20 208.889
R486 vdd.t20 vdd.t27 208.889
R487 vdd.t27 vdd.t14 208.889
R488 vdd.t14 vdd.t18 208.889
R489 vdd.t18 vdd.t25 208.889
R490 vdd.t25 vdd.t12 208.889
R491 vdd.t12 vdd.t21 208.889
R492 vdd.t21 vdd.t30 208.889
R493 vdd.t30 vdd.t15 208.889
R494 vdd.t15 vdd.t22 208.889
R495 vdd.n13 vdd.n8 13.3235
R496 vdd.n2 vdd.t6 9.66464
R497 vdd.n5 vdd.n1 6.96188
R498 vdd.n10 vdd.n9 6.29206
R499 vdd.n8 vdd.t8 5.27561
R500 vdd.n0 vdd.t4 5.26126
R501 vdd.n2 vdd.t11 3.69646
R502 vdd.n12 vdd.n11 3.54271
R503 vdd.n4 vdd.n3 3.13374
R504 vdd.n6 vdd.n0 2.43993
R505 vdd.n11 vdd.n7 2.08974
R506 vdd vdd.n14 1.83775
R507 vdd.n14 vdd.n13 1.61594
R508 vdd.n4 vdd.n2 1.60498
R509 vdd.n12 vdd.n10 0.698
R510 vdd.n13 vdd.n12 0.557375
R511 vdd.n5 vdd.n4 0.337689
R512 vdd.n6 vdd.n5 0.248933
R513 vdd.n14 vdd.n7 0.206214
R514 vdd.n7 vdd.n6 0.0067212
R515 clk.n3 clk.t0 35.7254
R516 clk.n0 clk.t6 35.7221
R517 clk.n2 clk.t3 34.0719
R518 clk.n4 clk.t2 30.1393
R519 clk.n1 clk.t5 30.1393
R520 clk.n5 clk.t1 26.8518
R521 clk.n3 clk.t4 15.823
R522 clk.n0 clk.t7 15.8225
R523 clk.n1 clk.n0 10.7103
R524 clk.n4 clk.n3 10.6727
R525 clk.n6 clk.n2 1.57407
R526 clk clk.n6 0.460065
R527 clk.n6 clk.n5 0.281711
R528 clk.n2 clk.n1 0.113703
R529 clk.n5 clk.n4 0.0995311
R530 nclk.n0 nclk.t7 35.0711
R531 nclk.n3 nclk.t1 28.37
R532 nclk.n1 nclk.t6 25.9811
R533 nclk.n3 nclk.t0 25.2836
R534 nclk.n5 nclk.t4 24.2876
R535 nclk.n2 nclk.t3 24.2876
R536 nclk.n4 nclk.t2 19.9399
R537 nclk.n0 nclk.t5 19.5588
R538 nclk.n2 nclk.n1 7.06888
R539 nclk.n5 nclk.n4 7.0647
R540 nclk.n6 nclk.n5 2.40549
R541 nclk.n6 nclk.n2 1.7803
R542 nclk.n4 nclk.n3 0.699125
R543 nclk nclk.n6 0.594832
R544 nclk.n1 nclk.n0 0.381269
C0 nclk a_5944_2919# 0.11947f
C1 vout vin 15.538f
C2 vdd a_5939_n1022# 0.47578f
C3 vin a_8039_2775# 0.50886f
C4 vout a_5939_n1022# 0.00174f
C5 vin a_8034_n1134# 0.23448f
C6 vout vdd 1.94458f
C7 vin clk 0.13055f
C8 vin nclk 1.44517f
C9 a_8034_n1134# a_5939_n1022# 0.91362f
C10 vdd a_8039_2775# 0.84309f
C11 vin a_5944_2919# 0.05645f
C12 vdd a_8034_n1134# 0.58164f
C13 clk a_5939_n1022# 0.99882f
C14 vout a_8039_2775# 0.00196f
C15 nclk a_5939_n1022# 0.12266f
C16 clk vdd 2.23886f
C17 nclk vdd 3.22814f
C18 vout a_8034_n1134# 0.00218f
C19 vdd a_5944_2919# 0.18588f
C20 vout clk 1.05144f
C21 vout nclk 0.17473f
C22 clk a_8039_2775# 0.68178f
C23 vout a_5944_2919# 0.00216f
C24 nclk a_8039_2775# 0.68724f
C25 a_8039_2775# a_5944_2919# 0.87176f
C26 clk a_8034_n1134# 0.65772f
C27 vin a_5939_n1022# 0.02754f
C28 nclk a_8034_n1134# 0.5632f
C29 vin vdd 1.55661f
C30 nclk clk 2.72524f
C31 clk a_5944_2919# 0.85419f
C32 vout vss 5.04024f
C33 vin vss 2.81869f
C34 nclk vss 6.76427f
C35 clk vss 8.52934f
C36 vdd vss 41.3125f
C37 a_8034_n1134# vss 4.44835f
C38 a_5939_n1022# vss 2.41334f
C39 a_8039_2775# vss 2.76621f
C40 a_5944_2919# vss 1.70938f
C41 nclk.t7 vss 0.02839f
C42 nclk.t5 vss 0.1214f
C43 nclk.n0 vss 0.25404f
C44 nclk.t6 vss 0.13476f
C45 nclk.n1 vss 0.48461f
C46 nclk.t3 vss 0.16661f
C47 nclk.n2 vss 0.58828f
C48 nclk.t2 vss 0.12284f
C49 nclk.t1 vss 0.02302f
C50 nclk.t0 vss 0.12928f
C51 nclk.n3 vss 0.48242f
C52 nclk.n4 vss 0.35941f
C53 nclk.t4 vss 0.16661f
C54 nclk.n5 vss 0.7867f
C55 nclk.n6 vss 1.61769f
C56 clk.t7 vss 0.04729f
C57 clk.t6 vss 0.13069f
C58 clk.n0 vss 0.31002f
C59 clk.t5 vss 0.14661f
C60 clk.n1 vss 0.44974f
C61 clk.t3 vss 0.01724f
C62 clk.n2 vss 0.83255f
C63 clk.t1 vss 0.00981f
C64 clk.t4 vss 0.04729f
C65 clk.t0 vss 0.13706f
C66 clk.n3 vss 0.31464f
C67 clk.t2 vss 0.14661f
C68 clk.n4 vss 0.45569f
C69 clk.n5 vss 0.3017f
C70 clk.n6 vss 1.17108f
C71 vdd.t4 vss 0.01071f
C72 vdd.n0 vss 0.09707f
C73 vdd.t3 vss 0.10128f
C74 vdd.n1 vss 0.12425f
C75 vdd.t6 vss 0.00937f
C76 vdd.t11 vss 0.01713f
C77 vdd.n2 vss 0.04998f
C78 vdd.t2 vss 0.17065f
C79 vdd.t10 vss 0.17147f
C80 vdd.t1 vss 0.17266f
C81 vdd.n3 vss 0.32172f
C82 vdd.n4 vss 0.09419f
C83 vdd.n5 vss 0.0972f
C84 vdd.n6 vss 0.07182f
C85 vdd.n7 vss 0.06243f
C86 vdd.t8 vss 0.01074f
C87 vdd.n8 vss 0.2186f
C88 vdd.t7 vss 0.12673f
C89 vdd.t0 vss 0.16408f
C90 vdd.n9 vss 0.3232f
C91 vdd.t9 vss 0.1708f
C92 vdd.t5 vss 0.17196f
C93 vdd.n10 vss 0.17072f
C94 vdd.t22 vss 0.20056f
C95 vdd.t15 vss 0.09333f
C96 vdd.t30 vss 0.09333f
C97 vdd.t21 vss 0.09333f
C98 vdd.t12 vss 0.09333f
C99 vdd.t25 vss 0.09333f
C100 vdd.t18 vss 0.09333f
C101 vdd.t14 vss 0.09333f
C102 vdd.t27 vss 0.09333f
C103 vdd.t20 vss 0.09333f
C104 vdd.t26 vss 0.09333f
C105 vdd.t19 vss 0.09333f
C106 vdd.t16 vss 0.09333f
C107 vdd.t29 vss 0.09333f
C108 vdd.t24 vss 0.09333f
C109 vdd.t13 vss 0.09333f
C110 vdd.t23 vss 0.09333f
C111 vdd.t17 vss 0.09333f
C112 vdd.t31 vss 0.09333f
C113 vdd.t28 vss 0.11513f
C114 vdd.n11 vss 0.19063f
C115 vdd.n12 vss 0.07661f
C116 vdd.n13 vss 2.13687f
C117 vdd.n14 vss 1.25285f
C118 a_5297_1329.n2 vss 0.0225f
C119 a_5297_1329.t13 vss 0.08905f
C120 a_5297_1329.t20 vss 0.08877f
C121 a_5297_1329.n3 vss 0.1212f
C122 a_5297_1329.t5 vss 0.08877f
C123 a_5297_1329.n4 vss 0.06522f
C124 a_5297_1329.t14 vss 0.08877f
C125 a_5297_1329.n5 vss 0.06522f
C126 a_5297_1329.t23 vss 0.08877f
C127 a_5297_1329.n6 vss 0.06522f
C128 a_5297_1329.t10 vss 0.08877f
C129 a_5297_1329.n7 vss 0.06522f
C130 a_5297_1329.t17 vss 0.08877f
C131 a_5297_1329.n8 vss 0.06522f
C132 a_5297_1329.t21 vss 0.08877f
C133 a_5297_1329.n9 vss 0.05775f
C134 a_5297_1329.n10 vss 0.02252f
C135 a_5297_1329.t15 vss 0.08877f
C136 a_5297_1329.n11 vss 0.05108f
C137 a_5297_1329.t8 vss 0.08877f
C138 a_5297_1329.n12 vss 0.05107f
C139 a_5297_1329.n13 vss 0.02251f
C140 a_5297_1329.t7 vss 0.08905f
C141 a_5297_1329.t4 vss 0.08877f
C142 a_5297_1329.n14 vss 0.1212f
C143 a_5297_1329.t18 vss 0.08877f
C144 a_5297_1329.n15 vss 0.06522f
C145 a_5297_1329.t12 vss 0.08877f
C146 a_5297_1329.n16 vss 0.06522f
C147 a_5297_1329.t22 vss 0.08877f
C148 a_5297_1329.n17 vss 0.06522f
C149 a_5297_1329.t11 vss 0.08877f
C150 a_5297_1329.n18 vss 0.06522f
C151 a_5297_1329.t6 vss 0.08877f
C152 a_5297_1329.n19 vss 0.06522f
C153 a_5297_1329.t19 vss 0.08877f
C154 a_5297_1329.n20 vss 0.06522f
C155 a_5297_1329.t16 vss 0.08877f
C156 a_5297_1329.n21 vss 0.0548f
C157 a_5297_1329.t9 vss 0.08877f
C158 a_5297_1329.n22 vss 0.0511f
C159 a_5297_1329.n23 vss 0.02246f
C160 a_5297_1329.n24 vss 0.82798f
C161 a_5297_1329.n25 vss 0.21069f
C162 a_5297_1329.t2 vss 0.0657f
C163 a_5297_1329.t1 vss 0.03559f
C164 a_5297_1329.n26 vss 0.15401f
C165 a_5297_1329.n27 vss 0.39189f
C166 a_5297_1329.n28 vss 0.21069f
C167 a_5297_1329.n29 vss 0.18815f
C168 a_5297_1329.n30 vss 0.89507f
C169 a_5297_1329.n31 vss 0.17358f
C170 a_5297_1329.t3 vss 0.03559f
C171 a_5297_1329.n32 vss 0.15383f
C172 a_5297_1329.t0 vss 0.06571f
C173 vout.n0 vss 0.11453f
C174 vout.t26 vss 0.27416f
C175 vout.t6 vss 0.22981f
C176 vout.n1 vss 0.71753f
C177 vout.t2 vss 0.04819f
C178 vout.t33 vss 0.04819f
C179 vout.n2 vss 0.1478f
C180 vout.t5 vss 0.04819f
C181 vout.t31 vss 0.04819f
C182 vout.n3 vss 0.1478f
C183 vout.t11 vss 0.06047f
C184 vout.t16 vss 0.06047f
C185 vout.n4 vss 0.18419f
C186 vout.n5 vss 0.33623f
C187 vout.n6 vss 0.11453f
C188 vout.t3 vss 0.04819f
C189 vout.t4 vss 0.04819f
C190 vout.n7 vss 0.1478f
C191 vout.t19 vss 0.06047f
C192 vout.t23 vss 0.06047f
C193 vout.n8 vss 0.18419f
C194 vout.n9 vss 0.11405f
C195 vout.n10 vss 0.11453f
C196 vout.t29 vss 0.04819f
C197 vout.t35 vss 0.04819f
C198 vout.n11 vss 0.1478f
C199 vout.t12 vss 0.06047f
C200 vout.t15 vss 0.06047f
C201 vout.n12 vss 0.18419f
C202 vout.t1 vss 0.04819f
C203 vout.t27 vss 0.04819f
C204 vout.n13 vss 0.1478f
C205 vout.t20 vss 0.06047f
C206 vout.t21 vss 0.06047f
C207 vout.n14 vss 0.18419f
C208 vout.n15 vss 0.33623f
C209 vout.n16 vss 0.11453f
C210 vout.t9 vss 0.04819f
C211 vout.t30 vss 0.04819f
C212 vout.n17 vss 0.1478f
C213 vout.t24 vss 0.06047f
C214 vout.t14 vss 0.06047f
C215 vout.n18 vss 0.18419f
C216 vout.n19 vss 0.11405f
C217 vout.n20 vss 0.11453f
C218 vout.t34 vss 0.04819f
C219 vout.t10 vss 0.04819f
C220 vout.n21 vss 0.1478f
C221 vout.t17 vss 0.06047f
C222 vout.t22 vss 0.06047f
C223 vout.n22 vss 0.18419f
C224 vout.t28 vss 0.04819f
C225 vout.t0 vss 0.04819f
C226 vout.n23 vss 0.1478f
C227 vout.t25 vss 0.06047f
C228 vout.t13 vss 0.06047f
C229 vout.n24 vss 0.18419f
C230 vout.n25 vss 0.33623f
C231 vout.n26 vss 0.20378f
C232 vout.t7 vss 0.04819f
C233 vout.t32 vss 0.04819f
C234 vout.n27 vss 0.1478f
C235 vout.t18 vss 0.27416f
C236 vout.t8 vss 0.22981f
C237 vout.n28 vss 0.7161f
C238 vout.n29 vss 0.01235f
C239 vout.n30 vss 0.18821f
C240 vout.n31 vss 0.10764f
C241 vout.n32 vss 0.0834f
C242 vout.n33 vss 0.11453f
C243 vout.n34 vss 0.11453f
C244 vout.n35 vss 0.08768f
C245 vout.n36 vss 0.10336f
C246 vout.n37 vss 0.33623f
C247 vout.n38 vss 0.06772f
C248 vout.n39 vss 0.11453f
C249 vout.n40 vss 0.11453f
C250 vout.n41 vss 0.11453f
C251 vout.n42 vss 0.06629f
C252 vout.n43 vss 0.33623f
C253 vout.n44 vss 0.10479f
C254 vout.n45 vss 0.08625f
C255 vout.n46 vss 0.11453f
C256 vout.n47 vss 0.11453f
C257 vout.n48 vss 0.08483f
C258 vout.n49 vss 0.10621f
C259 vout.n50 vss 0.33623f
C260 vout.n51 vss 0.06487f
C261 vout.n52 vss 0.11453f
C262 vout.n53 vss 0.11453f
C263 vout.n54 vss 0.11453f
C264 vout.n55 vss 0.06914f
C265 vout.n56 vss 0.33623f
C266 vout.n57 vss 0.10193f
C267 vout.n58 vss 0.0891f
C268 vout.n59 vss 0.11453f
C269 vout.n60 vss 0.11453f
C270 vout.n61 vss 0.08197f
C271 vout.n62 vss 0.10906f
C272 vout.n63 vss 0.18821f
C273 vout.n64 vss 0.00998f
C274 vout.n65 vss 1.03825f
C275 vin.n0 vss 0.56838f
C276 vin.t22 vss 0.03547f
C277 vin.t18 vss 0.03547f
C278 vin.n1 vss 0.11139f
C279 vin.n2 vss 0.20185f
C280 vin.t12 vss 0.02827f
C281 vin.t32 vss 0.02827f
C282 vin.n3 vss 0.08891f
C283 vin.n4 vss 0.09997f
C284 vin.n5 vss 0.56838f
C285 vin.t24 vss 0.03547f
C286 vin.t15 vss 0.03547f
C287 vin.n6 vss 0.11126f
C288 vin.n7 vss 0.13731f
C289 vin.n8 vss 0.56838f
C290 vin.t29 vss 0.02827f
C291 vin.t10 vss 0.02827f
C292 vin.n9 vss 0.08891f
C293 vin.n10 vss 0.09997f
C294 vin.n11 vss 0.56838f
C295 vin.t13 vss 0.03547f
C296 vin.t19 vss 0.03547f
C297 vin.n12 vss 0.11126f
C298 vin.n13 vss 0.13731f
C299 vin.n14 vss 0.56838f
C300 vin.t4 vss 0.02827f
C301 vin.t33 vss 0.02827f
C302 vin.n15 vss 0.08891f
C303 vin.n16 vss 0.09997f
C304 vin.n17 vss 0.56838f
C305 vin.n18 vss 0.11039f
C306 vin.n19 vss 0.56838f
C307 vin.t7 vss 0.02827f
C308 vin.t2 vss 0.02827f
C309 vin.n20 vss 0.09608f
C310 vin.t37 vss 0.02827f
C311 vin.t6 vss 0.02827f
C312 vin.n21 vss 0.08891f
C313 vin.n22 vss 0.43496f
C314 vin.n23 vss 0.10192f
C315 vin.t31 vss 0.042f
C316 vin.t5 vss 0.09045f
C317 vin.n24 vss 0.21223f
C318 vin.t30 vss 0.03103f
C319 vin.t11 vss 0.05022f
C320 vin.n25 vss 0.17269f
C321 vin.n26 vss 0.45112f
C322 vin.n27 vss 0.34437f
C323 vin.t27 vss 0.03547f
C324 vin.t16 vss 0.03547f
C325 vin.n28 vss 0.11185f
C326 vin.n29 vss 0.25268f
C327 vin.t20 vss 0.03547f
C328 vin.t25 vss 0.03547f
C329 vin.n30 vss 0.11126f
C330 vin.n31 vss 0.13731f
C331 vin.n32 vss 0.17395f
C332 vin.n33 vss 0.56838f
C333 vin.n34 vss 0.1359f
C334 vin.t35 vss 0.02827f
C335 vin.t3 vss 0.02827f
C336 vin.n35 vss 0.08891f
C337 vin.n36 vss 0.09997f
C338 vin.n37 vss 0.08624f
C339 vin.n38 vss 0.07753f
C340 vin.n39 vss 0.14809f
C341 vin.n40 vss 0.56838f
C342 vin.n41 vss 0.18956f
C343 vin.n42 vss 0.09924f
C344 vin.t26 vss 0.03547f
C345 vin.t14 vss 0.03547f
C346 vin.n43 vss 0.11126f
C347 vin.n44 vss 0.13731f
C348 vin.n45 vss 0.11931f
C349 vin.n46 vss 0.1851f
C350 vin.n47 vss 0.56838f
C351 vin.n48 vss 0.14461f
C352 vin.n49 vss 0.09321f
C353 vin.t39 vss 0.02827f
C354 vin.t1 vss 0.02827f
C355 vin.n50 vss 0.08891f
C356 vin.n51 vss 0.09997f
C357 vin.n52 vss 0.10889f
C358 vin.n53 vss 0.12893f
C359 vin.n54 vss 0.56838f
C360 vin.n55 vss 0.16503f
C361 vin.n56 vss 0.13938f
C362 vin.t17 vss 0.03547f
C363 vin.t28 vss 0.03547f
C364 vin.n57 vss 0.11126f
C365 vin.n58 vss 0.13731f
C366 vin.n59 vss 0.15945f
C367 vin.n60 vss 0.14496f
C368 vin.n61 vss 0.56838f
C369 vin.n62 vss 0.11325f
C370 vin.n63 vss 0.12457f
C371 vin.t34 vss 0.02827f
C372 vin.t38 vss 0.02827f
C373 vin.n64 vss 0.08891f
C374 vin.n65 vss 0.09997f
C375 vin.n66 vss 0.14025f
C376 vin.n67 vss 0.09757f
C377 vin.n68 vss 0.56838f
C378 vin.n69 vss 0.12489f
C379 vin.n70 vss 0.17952f
C380 vin.t21 vss 0.03547f
C381 vin.t23 vss 0.03547f
C382 vin.n71 vss 0.11126f
C383 vin.n72 vss 0.13731f
C384 vin.n73 vss 0.18956f
C385 vin.n74 vss 0.10482f
C386 vin.n75 vss 0.56838f
C387 vin.n76 vss 0.08189f
C388 vin.n77 vss 0.14809f
C389 vin.t36 vss 0.02827f
C390 vin.t9 vss 0.02827f
C391 vin.n78 vss 0.09608f
C392 vin.t0 vss 0.02827f
C393 vin.t8 vss 0.02827f
C394 vin.n79 vss 0.08891f
C395 vin.n80 vss 0.41492f
C396 vin.n81 vss 0.08189f
C397 vin.n82 vss 0.81513f
C398 a_5673_n171.n2 vss 0.07314f
C399 a_5673_n171.t3 vss 0.02281f
C400 a_5673_n171.t1 vss 0.01236f
C401 a_5673_n171.n3 vss 0.05347f
C402 a_5673_n171.n4 vss 0.00784f
C403 a_5673_n171.t12 vss 0.03818f
C404 a_5673_n171.t17 vss 0.03809f
C405 a_5673_n171.n5 vss 0.04758f
C406 a_5673_n171.t5 vss 0.03809f
C407 a_5673_n171.n6 vss 0.02544f
C408 a_5673_n171.t8 vss 0.03809f
C409 a_5673_n171.n7 vss 0.02544f
C410 a_5673_n171.t13 vss 0.03809f
C411 a_5673_n171.n8 vss 0.02544f
C412 a_5673_n171.t16 vss 0.03809f
C413 a_5673_n171.n9 vss 0.02272f
C414 a_5673_n171.n10 vss 0.00784f
C415 a_5673_n171.t9 vss 0.03809f
C416 a_5673_n171.n11 vss 0.02029f
C417 a_5673_n171.t6 vss 0.03809f
C418 a_5673_n171.n12 vss 0.02029f
C419 a_5673_n171.n13 vss 0.00784f
C420 a_5673_n171.t4 vss 0.03818f
C421 a_5673_n171.t19 vss 0.03809f
C422 a_5673_n171.n14 vss 0.04758f
C423 a_5673_n171.t14 vss 0.03809f
C424 a_5673_n171.n15 vss 0.02544f
C425 a_5673_n171.t11 vss 0.03809f
C426 a_5673_n171.n16 vss 0.02544f
C427 a_5673_n171.t7 vss 0.03809f
C428 a_5673_n171.n17 vss 0.02544f
C429 a_5673_n171.t18 vss 0.03809f
C430 a_5673_n171.n18 vss 0.02544f
C431 a_5673_n171.t15 vss 0.03809f
C432 a_5673_n171.n19 vss 0.02161f
C433 a_5673_n171.t10 vss 0.03809f
C434 a_5673_n171.n20 vss 0.02029f
C435 a_5673_n171.n21 vss 0.00784f
C436 a_5673_n171.n22 vss 0.26925f
C437 a_5673_n171.n23 vss 0.29043f
C438 a_5673_n171.n24 vss 0.07314f
C439 a_5673_n171.n25 vss 0.06532f
C440 a_5673_n171.n26 vss 0.07178f
C441 a_5673_n171.n27 vss 0.06026f
C442 a_5673_n171.t2 vss 0.01236f
C443 a_5673_n171.n28 vss 0.0534f
C444 a_5673_n171.t0 vss 0.02281f
.ends

